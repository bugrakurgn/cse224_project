* NGSPICE file created from alu.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

.subckt alu VGND VPWR din1[0] din1[1] din1[2] din1[3] din1[4] din1[5] din1[6] din1[7]
+ din2[0] din2[1] din2[2] din2[3] din2[4] din2[5] din2[6] din2[7] dout[0] dout[1]
+ dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] op[0] op[1] op[2]
XFILLER_0_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_294_ _048_ _049_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_15_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_346_ _089_ _092_ _096_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__or3_4
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_277_ _033_ _023_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__and2b_1
X_200_ _117_ _127_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__nand2_1
X_329_ _079_ _080_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput20 net20 VGND VGND VPWR VPWR dout[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_18_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_293_ net15 _025_ net28 VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_21_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_276_ _019_ _166_ _015_ _030_ _029_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__a311oi_4
X_345_ _138_ _100_ _093_ _095_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_328_ _169_ _008_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__nand2_1
X_259_ net14 _016_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_24_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput21 net21 VGND VGND VPWR VPWR dout[1] sky130_fd_sc_hd__buf_2
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_292_ net16 net8 VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__xnor2_2
X_344_ net13 net5 _094_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__a21oi_1
X_275_ _029_ _031_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_189_ _102_ _116_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__xnor2_4
X_258_ net13 net28 _164_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__a21o_1
X_327_ _012_ _011_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput22 net22 VGND VGND VPWR VPWR dout[2] sky130_fd_sc_hd__buf_2
XFILLER_0_27_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_291_ _032_ _034_ _047_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__a21o_1
XFILLER_0_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_274_ _019_ _166_ _015_ _030_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__a31o_1
X_343_ net5 _153_ _090_ _158_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_257_ _008_ _169_ _011_ _012_ _014_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__a311o_4
X_326_ _008_ _023_ _072_ _078_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__a31o_1
X_188_ _110_ _115_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_9_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_309_ _101_ _103_ _156_ _062_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput23 net23 VGND VGND VPWR VPWR dout[3] sky130_fd_sc_hd__buf_2
XFILLER_0_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_290_ _100_ _040_ _041_ _046_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_273_ _018_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__inv_2
X_342_ _134_ _137_ _129_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_187_ _111_ _113_ _114_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__o21bai_4
X_256_ _166_ _013_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _134_ _073_ _077_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__o21bai_2
X_239_ _163_ _162_ _106_ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_308_ _101_ _103_ _158_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_10_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput24 net24 VGND VGND VPWR VPWR dout[4] sky130_fd_sc_hd__buf_2
XFILLER_0_12_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_341_ net13 net5 _151_ _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__a31o_1
X_272_ _027_ _028_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_0_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_255_ net5 _165_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__or2_1
X_186_ net9 net10 net3 net4 VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__and4_1
X_324_ _104_ _106_ _151_ _075_ _076_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__a311o_1
XFILLER_0_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_307_ _112_ _118_ _058_ _061_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__a31o_1
XFILLER_0_21_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_238_ net5 _165_ VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__nand2_2
XFILLER_0_1_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput25 net25 VGND VGND VPWR VPWR dout[5] sky130_fd_sc_hd__buf_2
XFILLER_0_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_340_ _090_ _156_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_271_ net7 _026_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_254_ _107_ _010_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__nor2_1
X_323_ _104_ _153_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__nor2_1
X_185_ _103_ net3 net4 _112_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_237_ net13 _164_ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_306_ _118_ _153_ _060_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput26 net26 VGND VGND VPWR VPWR dout[6] sky130_fd_sc_hd__buf_2
XFILLER_0_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_270_ net7 _026_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_322_ _104_ _106_ _156_ _074_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__o22a_1
X_184_ net9 VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_253_ _107_ _010_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_305_ _112_ _118_ _155_ _059_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__a31o_1
X_236_ net11 net12 _162_ _163_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__o31a_2
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_219_ _128_ _138_ _146_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__a21oi_1
Xoutput27 net27 VGND VGND VPWR VPWR dout[7] sky130_fd_sc_hd__buf_2
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_252_ _119_ _009_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__xnor2_2
X_321_ _104_ _106_ _158_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__a21oi_1
X_183_ net2 net11 VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_235_ net17 net18 net19 VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_18_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_304_ _112_ _118_ _099_ _150_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_218_ _144_ _145_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__or2b_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_320_ _132_ _133_ _100_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__o21ai_2
X_182_ _105_ _108_ _109_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__o21ai_4
X_251_ _106_ _162_ net28 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_303_ _100_ _151_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_23_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_234_ net9 net10 VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__or2_4
XFILLER_0_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_217_ _139_ _140_ _143_ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_181_ _104_ _106_ net4 _103_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__a22o_1
X_250_ _002_ _005_ _007_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_302_ _023_ _051_ _052_ _057_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__a31o_1
X_233_ net14 net6 _151_ _154_ _160_ VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__a311o_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_216_ _139_ _140_ _143_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__nor3_1
XFILLER_0_20_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_180_ _106_ _107_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__nand2_2
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_232_ net14 net6 _156_ _159_ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__o22a_1
X_301_ _100_ _053_ _056_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_215_ _141_ _142_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_6_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_300_ net8 _153_ _048_ _158_ _055_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__o221a_1
X_231_ net14 net6 _158_ VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__a21oi_1
Xinput1 din1[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_27_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_214_ _104_ _119_ VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_6_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_230_ _157_ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__buf_2
XFILLER_0_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 din1[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
X_213_ _106_ _107_ _105_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_2_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 din1[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_289_ net7 _153_ _044_ _045_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__o211ai_1
X_212_ _101_ _119_ _116_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 din1[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
X_288_ net18 _043_ _042_ _155_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_211_ _110_ _115_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_287_ _158_ _042_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__or3b_1
Xinput5 din1[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
X_210_ _129_ _134_ _137_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__nand3_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_339_ net13 net5 VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_286_ net15 net7 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 din1[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_269_ net15 _025_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__xnor2_1
X_338_ _015_ _023_ _088_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_285_ net15 net7 VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 din1[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_268_ net14 net13 _164_ net28 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__o31a_1
X_199_ _118_ _119_ _125_ _126_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__a31o_1
X_337_ _014_ _087_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput10 din2[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_22_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_284_ _038_ _039_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 din1[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_198_ _120_ _121_ _124_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__and3_1
X_267_ _100_ _149_ _161_ _024_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__a211o_1
X_336_ _169_ _008_ _011_ _012_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_319_ _007_ _002_ _005_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__or3_1
Xinput11 din2[2] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 din2[0] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_1_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _038_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_197_ _120_ _121_ _124_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_266_ _021_ _022_ _023_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__and3_1
X_335_ _023_ _081_ _082_ _100_ _086_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__a221o_1
XFILLER_0_2_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 din2[3] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
X_249_ _169_ _006_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__and2_2
X_318_ _071_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_282_ _128_ _145_ _144_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_334_ _119_ _107_ _151_ _084_ _085_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__a311o_1
X_196_ net1 _106_ _122_ _123_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__a31o_1
X_265_ net19 _099_ _150_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__and3_2
XFILLER_0_2_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_179_ net4 VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__clkbuf_4
Xinput13 din2[4] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_317_ _063_ _066_ _067_ _070_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_248_ _104_ _167_ _168_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_281_ _036_ _037_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_264_ _020_ _166_ _015_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__nand3_1
X_333_ _107_ _153_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_195_ net9 net2 net10 net3 VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_316_ _005_ _069_ _023_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__or3b_1
Xinput14 din2[5] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
X_247_ _002_ _003_ _004_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__and3b_2
X_178_ net11 VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_280_ _119_ _107_ _035_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_332_ _119_ _107_ _156_ _083_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_194_ net2 net10 _104_ _112_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__a22o_1
X_263_ _166_ _015_ _020_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput15 din2[6] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
X_177_ _103_ _104_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__nand2_2
X_315_ _068_ _004_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__nor2_1
X_246_ _118_ _112_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_229_ net17 net19 net18 VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_262_ _018_ _019_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__nand2_1
X_331_ _119_ _107_ _158_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__a21oi_1
X_193_ _114_ _113_ _111_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_245_ _101_ _000_ _001_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__or3_4
X_176_ net3 VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__buf_4
Xinput16 din2[7] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
X_314_ _002_ _003_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_228_ net18 _155_ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__nor2_2
XFILLER_0_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone1 net17 net18 net19 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__nand3b_2
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_330_ _134_ _137_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__xor2_1
X_192_ _114_ _111_ _113_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__or3_1
X_261_ net6 _017_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_244_ _000_ _001_ _101_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__o21a_2
X_175_ net10 VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_16_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_313_ _101_ _153_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nor2_1
Xinput17 op[0] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_227_ net17 _098_ VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__nand2_2
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_260_ net6 _017_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_191_ net12 VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_243_ _112_ _163_ _103_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__a21oi_1
X_312_ _101_ _103_ _151_ _065_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_16_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 op[1] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_4
X_174_ _101_ net12 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__nand2_2
XFILLER_0_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_226_ net6 _153_ VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_209_ _135_ _136_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_190_ net1 VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 op[2] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_4
X_311_ _133_ _100_ _064_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__and3b_1
XFILLER_0_5_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_173_ net2 VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__clkbuf_4
X_242_ _112_ _103_ _163_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_225_ _152_ VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_9_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_208_ _126_ _125_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _112_ _101_ _103_ _118_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__a22o_1
X_241_ _167_ _168_ _104_ VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__o21ai_4
X_172_ _098_ _099_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_21_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_224_ net19 _099_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_25_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_207_ _118_ _119_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_171_ net17 net18 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__or2_2
X_240_ net11 _163_ _162_ VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_223_ net19 _150_ VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__nor2_4
XFILLER_0_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_206_ _132_ _133_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__and2_2
XFILLER_0_9_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ net19 VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_299_ net16 net8 _151_ _054_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__a31oi_1
X_222_ net17 net18 VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_205_ _112_ _118_ _101_ _103_ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_298_ net16 net8 _156_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_221_ _147_ _148_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_204_ _130_ _131_ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 _069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_297_ _038_ _039_ _036_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_220_ _128_ _138_ _146_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_8_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_203_ _123_ _122_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_2 _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_296_ _027_ _033_ _050_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_15_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_279_ _119_ _107_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nand3_1
X_202_ _118_ _106_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_295_ _027_ _033_ _050_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_12_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_278_ _105_ _142_ _108_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_347_ _097_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
X_201_ _117_ _127_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

