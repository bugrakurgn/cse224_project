VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu
  CLASS BLOCK ;
  FOREIGN alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.020 10.640 39.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.020 10.640 64.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.020 10.640 89.620 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.380 94.540 19.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 43.380 94.540 44.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 68.380 94.540 69.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.720 10.640 36.320 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.720 10.640 61.320 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.720 10.640 86.320 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.080 94.540 16.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 40.080 94.540 41.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 65.080 94.540 66.680 ;
    END
  END VPWR
  PIN din1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END din1[0]
  PIN din1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END din1[1]
  PIN din1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END din1[2]
  PIN din1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END din1[3]
  PIN din1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END din1[4]
  PIN din1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END din1[5]
  PIN din1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END din1[6]
  PIN din1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END din1[7]
  PIN din2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END din2[0]
  PIN din2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END din2[1]
  PIN din2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END din2[2]
  PIN din2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END din2[3]
  PIN din2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END din2[4]
  PIN din2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END din2[5]
  PIN din2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END din2[6]
  PIN din2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END din2[7]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 92.520 100.000 93.120 ;
    END
  END dout[0]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 80.280 100.000 80.880 ;
    END
  END dout[1]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 68.040 100.000 68.640 ;
    END
  END dout[2]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.800 100.000 56.400 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 43.560 100.000 44.160 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 31.320 100.000 31.920 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 19.080 100.000 19.680 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 6.840 100.000 7.440 ;
    END
  END dout[7]
  PIN op[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END op[0]
  PIN op[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END op[1]
  PIN op[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END op[2]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 94.490 87.125 ;
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 4.210 10.640 95.150 88.360 ;
      LAYER met2 ;
        RECT 4.230 4.280 95.120 93.005 ;
        RECT 4.230 4.000 16.370 4.280 ;
        RECT 17.210 4.000 49.490 4.280 ;
        RECT 50.330 4.000 82.610 4.280 ;
        RECT 83.450 4.000 95.120 4.280 ;
      LAYER met3 ;
        RECT 3.990 92.120 95.600 92.985 ;
        RECT 3.990 90.800 96.000 92.120 ;
        RECT 4.400 89.400 96.000 90.800 ;
        RECT 3.990 85.360 96.000 89.400 ;
        RECT 4.400 83.960 96.000 85.360 ;
        RECT 3.990 81.280 96.000 83.960 ;
        RECT 3.990 79.920 95.600 81.280 ;
        RECT 4.400 79.880 95.600 79.920 ;
        RECT 4.400 78.520 96.000 79.880 ;
        RECT 3.990 74.480 96.000 78.520 ;
        RECT 4.400 73.080 96.000 74.480 ;
        RECT 3.990 69.040 96.000 73.080 ;
        RECT 4.400 67.640 95.600 69.040 ;
        RECT 3.990 63.600 96.000 67.640 ;
        RECT 4.400 62.200 96.000 63.600 ;
        RECT 3.990 58.160 96.000 62.200 ;
        RECT 4.400 56.800 96.000 58.160 ;
        RECT 4.400 56.760 95.600 56.800 ;
        RECT 3.990 55.400 95.600 56.760 ;
        RECT 3.990 52.720 96.000 55.400 ;
        RECT 4.400 51.320 96.000 52.720 ;
        RECT 3.990 47.280 96.000 51.320 ;
        RECT 4.400 45.880 96.000 47.280 ;
        RECT 3.990 44.560 96.000 45.880 ;
        RECT 3.990 43.160 95.600 44.560 ;
        RECT 3.990 41.840 96.000 43.160 ;
        RECT 4.400 40.440 96.000 41.840 ;
        RECT 3.990 36.400 96.000 40.440 ;
        RECT 4.400 35.000 96.000 36.400 ;
        RECT 3.990 32.320 96.000 35.000 ;
        RECT 3.990 30.960 95.600 32.320 ;
        RECT 4.400 30.920 95.600 30.960 ;
        RECT 4.400 29.560 96.000 30.920 ;
        RECT 3.990 25.520 96.000 29.560 ;
        RECT 4.400 24.120 96.000 25.520 ;
        RECT 3.990 20.080 96.000 24.120 ;
        RECT 4.400 18.680 95.600 20.080 ;
        RECT 3.990 14.640 96.000 18.680 ;
        RECT 4.400 13.240 96.000 14.640 ;
        RECT 3.990 9.200 96.000 13.240 ;
        RECT 4.400 7.840 96.000 9.200 ;
        RECT 4.400 7.800 95.600 7.840 ;
        RECT 3.990 6.975 95.600 7.800 ;
      LAYER met4 ;
        RECT 12.255 11.735 12.620 85.505 ;
        RECT 15.020 11.735 34.320 85.505 ;
        RECT 36.720 11.735 37.620 85.505 ;
        RECT 40.020 11.735 59.320 85.505 ;
        RECT 61.720 11.735 62.620 85.505 ;
        RECT 65.020 11.735 84.320 85.505 ;
        RECT 86.720 11.735 87.105 85.505 ;
  END
END alu
END LIBRARY

