magic
tech sky130A
magscale 1 2
timestamp 1746363044
<< nwell >>
rect 1066 2159 18898 17425
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 842 2128 19030 17672
<< metal2 >>
rect 3330 0 3386 800
rect 9954 0 10010 800
rect 16578 0 16634 800
<< obsm2 >>
rect 846 856 19024 18601
rect 846 800 3274 856
rect 3442 800 9898 856
rect 10066 800 16522 856
rect 16690 800 19024 856
<< metal3 >>
rect 19200 18504 20000 18624
rect 0 17960 800 18080
rect 0 16872 800 16992
rect 19200 16056 20000 16176
rect 0 15784 800 15904
rect 0 14696 800 14816
rect 0 13608 800 13728
rect 19200 13608 20000 13728
rect 0 12520 800 12640
rect 0 11432 800 11552
rect 19200 11160 20000 11280
rect 0 10344 800 10464
rect 0 9256 800 9376
rect 19200 8712 20000 8832
rect 0 8168 800 8288
rect 0 7080 800 7200
rect 19200 6264 20000 6384
rect 0 5992 800 6112
rect 0 4904 800 5024
rect 0 3816 800 3936
rect 19200 3816 20000 3936
rect 0 2728 800 2848
rect 0 1640 800 1760
rect 19200 1368 20000 1488
<< obsm3 >>
rect 798 18424 19120 18597
rect 798 18160 19200 18424
rect 880 17880 19200 18160
rect 798 17072 19200 17880
rect 880 16792 19200 17072
rect 798 16256 19200 16792
rect 798 15984 19120 16256
rect 880 15976 19120 15984
rect 880 15704 19200 15976
rect 798 14896 19200 15704
rect 880 14616 19200 14896
rect 798 13808 19200 14616
rect 880 13528 19120 13808
rect 798 12720 19200 13528
rect 880 12440 19200 12720
rect 798 11632 19200 12440
rect 880 11360 19200 11632
rect 880 11352 19120 11360
rect 798 11080 19120 11352
rect 798 10544 19200 11080
rect 880 10264 19200 10544
rect 798 9456 19200 10264
rect 880 9176 19200 9456
rect 798 8912 19200 9176
rect 798 8632 19120 8912
rect 798 8368 19200 8632
rect 880 8088 19200 8368
rect 798 7280 19200 8088
rect 880 7000 19200 7280
rect 798 6464 19200 7000
rect 798 6192 19120 6464
rect 880 6184 19120 6192
rect 880 5912 19200 6184
rect 798 5104 19200 5912
rect 880 4824 19200 5104
rect 798 4016 19200 4824
rect 880 3736 19120 4016
rect 798 2928 19200 3736
rect 880 2648 19200 2928
rect 798 1840 19200 2648
rect 880 1568 19200 1840
rect 880 1560 19120 1568
rect 798 1395 19120 1560
<< metal4 >>
rect 1944 2128 2264 17456
rect 2604 2128 2924 17456
rect 6944 2128 7264 17456
rect 7604 2128 7924 17456
rect 11944 2128 12264 17456
rect 12604 2128 12924 17456
rect 16944 2128 17264 17456
rect 17604 2128 17924 17456
<< obsm4 >>
rect 2451 2347 2524 17101
rect 3004 2347 6864 17101
rect 7344 2347 7524 17101
rect 8004 2347 11864 17101
rect 12344 2347 12524 17101
rect 13004 2347 16864 17101
rect 17344 2347 17421 17101
<< metal5 >>
rect 1056 13676 18908 13996
rect 1056 13016 18908 13336
rect 1056 8676 18908 8996
rect 1056 8016 18908 8336
rect 1056 3676 18908 3996
rect 1056 3016 18908 3336
<< labels >>
rlabel metal4 s 2604 2128 2924 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17604 2128 17924 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3676 18908 3996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8676 18908 8996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 13676 18908 13996 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16944 2128 17264 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3016 18908 3336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8016 18908 8336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 13016 18908 13336 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 9256 800 9376 6 din1[0]
port 3 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 din1[1]
port 4 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 din1[2]
port 5 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 din1[3]
port 6 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 din1[4]
port 7 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 din1[5]
port 8 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 din1[6]
port 9 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 din1[7]
port 10 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 din2[0]
port 11 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 din2[1]
port 12 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 din2[2]
port 13 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 din2[3]
port 14 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 din2[4]
port 15 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 din2[5]
port 16 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 din2[6]
port 17 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 din2[7]
port 18 nsew signal input
rlabel metal3 s 19200 18504 20000 18624 6 dout[0]
port 19 nsew signal output
rlabel metal3 s 19200 16056 20000 16176 6 dout[1]
port 20 nsew signal output
rlabel metal3 s 19200 13608 20000 13728 6 dout[2]
port 21 nsew signal output
rlabel metal3 s 19200 11160 20000 11280 6 dout[3]
port 22 nsew signal output
rlabel metal3 s 19200 8712 20000 8832 6 dout[4]
port 23 nsew signal output
rlabel metal3 s 19200 6264 20000 6384 6 dout[5]
port 24 nsew signal output
rlabel metal3 s 19200 3816 20000 3936 6 dout[6]
port 25 nsew signal output
rlabel metal3 s 19200 1368 20000 1488 6 dout[7]
port 26 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 op[0]
port 27 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 op[1]
port 28 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 op[2]
port 29 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1279828
string GDS_FILE /openlane/designs/alu/runs/RUN_2025.05.04_12.49.18/results/signoff/alu.magic.gds
string GDS_START 434896
<< end >>

