magic
tech sky130A
magscale 1 2
timestamp 1746363043
<< viali >>
rect 18429 17289 18463 17323
rect 1869 17221 1903 17255
rect 2881 17221 2915 17255
rect 1501 17153 1535 17187
rect 2513 17153 2547 17187
rect 2789 17153 2823 17187
rect 5365 17153 5399 17187
rect 14749 17153 14783 17187
rect 15577 17153 15611 17187
rect 18245 17153 18279 17187
rect 15209 17085 15243 17119
rect 16037 17085 16071 17119
rect 1685 17017 1719 17051
rect 1961 16949 1995 16983
rect 5273 16949 5307 16983
rect 5549 16745 5583 16779
rect 15669 16745 15703 16779
rect 18153 16745 18187 16779
rect 4169 16677 4203 16711
rect 9965 16677 9999 16711
rect 10609 16677 10643 16711
rect 14933 16677 14967 16711
rect 6653 16609 6687 16643
rect 6837 16609 6871 16643
rect 6929 16609 6963 16643
rect 13553 16609 13587 16643
rect 14105 16609 14139 16643
rect 14657 16609 14691 16643
rect 15761 16609 15795 16643
rect 17049 16609 17083 16643
rect 5549 16541 5583 16575
rect 5733 16541 5767 16575
rect 6745 16541 6779 16575
rect 8493 16541 8527 16575
rect 8953 16541 8987 16575
rect 9137 16541 9171 16575
rect 9689 16541 9723 16575
rect 10333 16541 10367 16575
rect 12817 16541 12851 16575
rect 13093 16541 13127 16575
rect 14473 16541 14507 16575
rect 14749 16541 14783 16575
rect 14933 16541 14967 16575
rect 15025 16541 15059 16575
rect 15209 16541 15243 16575
rect 15669 16541 15703 16575
rect 16497 16541 16531 16575
rect 16589 16541 16623 16575
rect 16773 16541 16807 16575
rect 16865 16541 16899 16575
rect 17601 16541 17635 16575
rect 3801 16473 3835 16507
rect 7481 16473 7515 16507
rect 9965 16473 9999 16507
rect 10609 16473 10643 16507
rect 14197 16473 14231 16507
rect 15117 16473 15151 16507
rect 18337 16473 18371 16507
rect 4261 16405 4295 16439
rect 7113 16405 7147 16439
rect 9045 16405 9079 16439
rect 9781 16405 9815 16439
rect 10425 16405 10459 16439
rect 16037 16405 16071 16439
rect 17785 16405 17819 16439
rect 17969 16405 18003 16439
rect 18137 16405 18171 16439
rect 1685 16201 1719 16235
rect 17877 16201 17911 16235
rect 1961 16133 1995 16167
rect 12817 16133 12851 16167
rect 1501 16065 1535 16099
rect 1777 16065 1811 16099
rect 3065 16065 3099 16099
rect 3525 16065 3559 16099
rect 9597 16065 9631 16099
rect 11805 16065 11839 16099
rect 11897 16065 11931 16099
rect 13185 16065 13219 16099
rect 13369 16065 13403 16099
rect 13553 16065 13587 16099
rect 17785 16065 17819 16099
rect 18245 16065 18279 16099
rect 4353 15997 4387 16031
rect 9413 15997 9447 16031
rect 9505 15997 9539 16031
rect 9689 15997 9723 16031
rect 12081 15997 12115 16031
rect 1501 15929 1535 15963
rect 2145 15929 2179 15963
rect 9873 15861 9907 15895
rect 12265 15861 12299 15895
rect 13461 15861 13495 15895
rect 14197 15657 14231 15691
rect 14933 15657 14967 15691
rect 10517 15521 10551 15555
rect 10977 15521 11011 15555
rect 13553 15521 13587 15555
rect 17325 15521 17359 15555
rect 18429 15521 18463 15555
rect 6653 15453 6687 15487
rect 6745 15453 6779 15487
rect 8125 15453 8159 15487
rect 8309 15453 8343 15487
rect 10609 15453 10643 15487
rect 14105 15453 14139 15487
rect 14473 15453 14507 15487
rect 15485 15453 15519 15487
rect 16773 15453 16807 15487
rect 17141 15453 17175 15487
rect 17969 15453 18003 15487
rect 18245 15453 18279 15487
rect 13001 15385 13035 15419
rect 15117 15385 15151 15419
rect 15301 15385 15335 15419
rect 16865 15385 16899 15419
rect 6101 15317 6135 15351
rect 8217 15317 8251 15351
rect 14657 15317 14691 15351
rect 18061 15317 18095 15351
rect 8217 15113 8251 15147
rect 1501 14977 1535 15011
rect 3341 14977 3375 15011
rect 3525 14977 3559 15011
rect 5641 14977 5675 15011
rect 5733 14977 5767 15011
rect 7665 14977 7699 15011
rect 7941 14977 7975 15011
rect 8125 14977 8159 15011
rect 8309 14977 8343 15011
rect 9689 14977 9723 15011
rect 9965 14977 9999 15011
rect 13369 14977 13403 15011
rect 13921 14977 13955 15011
rect 14473 14977 14507 15011
rect 16865 14977 16899 15011
rect 16957 14977 16991 15011
rect 17233 14977 17267 15011
rect 9413 14909 9447 14943
rect 9873 14909 9907 14943
rect 10057 14909 10091 14943
rect 10148 14909 10182 14943
rect 15209 14909 15243 14943
rect 1685 14841 1719 14875
rect 7757 14841 7791 14875
rect 7849 14841 7883 14875
rect 9137 14841 9171 14875
rect 14841 14841 14875 14875
rect 3249 14773 3283 14807
rect 5917 14773 5951 14807
rect 7481 14773 7515 14807
rect 9505 14773 9539 14807
rect 10333 14773 10367 14807
rect 13737 14773 13771 14807
rect 14749 14773 14783 14807
rect 16681 14773 16715 14807
rect 17141 14773 17175 14807
rect 10149 14569 10183 14603
rect 9413 14501 9447 14535
rect 16681 14501 16715 14535
rect 10333 14433 10367 14467
rect 10057 14365 10091 14399
rect 14657 14365 14691 14399
rect 14841 14365 14875 14399
rect 16865 14365 16899 14399
rect 17141 14365 17175 14399
rect 9137 14297 9171 14331
rect 10333 14297 10367 14331
rect 9597 14229 9631 14263
rect 15669 14229 15703 14263
rect 17049 14229 17083 14263
rect 9229 14025 9263 14059
rect 18429 14025 18463 14059
rect 12449 13957 12483 13991
rect 12633 13957 12667 13991
rect 1409 13889 1443 13923
rect 8769 13889 8803 13923
rect 9045 13889 9079 13923
rect 13921 13889 13955 13923
rect 14565 13889 14599 13923
rect 14657 13889 14691 13923
rect 14841 13889 14875 13923
rect 18245 13889 18279 13923
rect 8861 13821 8895 13855
rect 8953 13821 8987 13855
rect 13645 13821 13679 13855
rect 13829 13821 13863 13855
rect 15025 13753 15059 13787
rect 1593 13685 1627 13719
rect 12265 13685 12299 13719
rect 13921 13685 13955 13719
rect 9045 13481 9079 13515
rect 13185 13481 13219 13515
rect 9325 13413 9359 13447
rect 9413 13413 9447 13447
rect 6929 13345 6963 13379
rect 12817 13345 12851 13379
rect 13001 13345 13035 13379
rect 14749 13345 14783 13379
rect 15945 13345 15979 13379
rect 3157 13277 3191 13311
rect 3341 13277 3375 13311
rect 3525 13277 3559 13311
rect 7021 13277 7055 13311
rect 9229 13277 9263 13311
rect 9505 13277 9539 13311
rect 12725 13277 12759 13311
rect 12909 13277 12943 13311
rect 14565 13277 14599 13311
rect 15485 13277 15519 13311
rect 15577 13277 15611 13311
rect 15117 13209 15151 13243
rect 1593 12937 1627 12971
rect 3065 12937 3099 12971
rect 7389 12937 7423 12971
rect 10517 12937 10551 12971
rect 6101 12869 6135 12903
rect 1409 12801 1443 12835
rect 3341 12801 3375 12835
rect 3801 12801 3835 12835
rect 4169 12801 4203 12835
rect 4537 12801 4571 12835
rect 4905 12801 4939 12835
rect 5457 12801 5491 12835
rect 5733 12801 5767 12835
rect 7021 12801 7055 12835
rect 7297 12801 7331 12835
rect 7757 12801 7791 12835
rect 8125 12801 8159 12835
rect 8309 12801 8343 12835
rect 10425 12801 10459 12835
rect 10517 12801 10551 12835
rect 13737 12801 13771 12835
rect 13829 12801 13863 12835
rect 6837 12733 6871 12767
rect 7665 12733 7699 12767
rect 13645 12733 13679 12767
rect 13921 12733 13955 12767
rect 7205 12665 7239 12699
rect 7757 12597 7791 12631
rect 8217 12597 8251 12631
rect 13461 12597 13495 12631
rect 9597 12393 9631 12427
rect 15117 12393 15151 12427
rect 7573 12325 7607 12359
rect 14657 12325 14691 12359
rect 9689 12257 9723 12291
rect 13369 12257 13403 12291
rect 14197 12257 14231 12291
rect 14381 12257 14415 12291
rect 2237 12189 2271 12223
rect 7113 12189 7147 12223
rect 7297 12189 7331 12223
rect 7757 12189 7791 12223
rect 8217 12189 8251 12223
rect 8309 12189 8343 12223
rect 8493 12189 8527 12223
rect 9413 12189 9447 12223
rect 9505 12189 9539 12223
rect 10333 12189 10367 12223
rect 11529 12189 11563 12223
rect 11713 12189 11747 12223
rect 11805 12189 11839 12223
rect 12173 12189 12207 12223
rect 13001 12189 13035 12223
rect 13185 12183 13219 12217
rect 13277 12189 13311 12223
rect 13553 12189 13587 12223
rect 14289 12189 14323 12223
rect 14473 12189 14507 12223
rect 15209 12189 15243 12223
rect 10149 12121 10183 12155
rect 10701 12121 10735 12155
rect 13737 12121 13771 12155
rect 2329 12053 2363 12087
rect 7113 12053 7147 12087
rect 8677 12053 8711 12087
rect 14749 12053 14783 12087
rect 11989 11781 12023 11815
rect 14289 11781 14323 11815
rect 1501 11713 1535 11747
rect 3893 11713 3927 11747
rect 3985 11713 4019 11747
rect 7205 11713 7239 11747
rect 7297 11713 7331 11747
rect 7481 11713 7515 11747
rect 10333 11713 10367 11747
rect 12173 11713 12207 11747
rect 14473 11713 14507 11747
rect 14657 11713 14691 11747
rect 17785 11713 17819 11747
rect 18245 11713 18279 11747
rect 10241 11645 10275 11679
rect 17509 11645 17543 11679
rect 17601 11645 17635 11679
rect 17693 11645 17727 11679
rect 1685 11577 1719 11611
rect 17969 11577 18003 11611
rect 3985 11509 4019 11543
rect 7665 11509 7699 11543
rect 10057 11509 10091 11543
rect 11805 11509 11839 11543
rect 18429 11509 18463 11543
rect 5917 11305 5951 11339
rect 15301 11305 15335 11339
rect 16037 11237 16071 11271
rect 2145 11169 2179 11203
rect 12541 11169 12575 11203
rect 14105 11169 14139 11203
rect 14289 11169 14323 11203
rect 14473 11169 14507 11203
rect 14841 11169 14875 11203
rect 14933 11169 14967 11203
rect 15025 11169 15059 11203
rect 15117 11169 15151 11203
rect 2329 11101 2363 11135
rect 2513 11101 2547 11135
rect 2605 11101 2639 11135
rect 4445 11101 4479 11135
rect 4813 11101 4847 11135
rect 5089 11101 5123 11135
rect 5917 11101 5951 11135
rect 6009 11101 6043 11135
rect 12265 11101 12299 11135
rect 12357 11101 12391 11135
rect 14381 11101 14415 11135
rect 14565 11101 14599 11135
rect 16221 11101 16255 11135
rect 5365 11033 5399 11067
rect 15945 11033 15979 11067
rect 16129 11033 16163 11067
rect 6285 10965 6319 10999
rect 12541 10965 12575 10999
rect 4077 10761 4111 10795
rect 4721 10761 4755 10795
rect 4997 10761 5031 10795
rect 1501 10693 1535 10727
rect 3801 10693 3835 10727
rect 4353 10693 4387 10727
rect 4813 10693 4847 10727
rect 1685 10625 1719 10659
rect 1777 10625 1811 10659
rect 1961 10625 1995 10659
rect 3985 10625 4019 10659
rect 4077 10625 4111 10659
rect 4169 10625 4203 10659
rect 4445 10625 4479 10659
rect 4537 10625 4571 10659
rect 5273 10625 5307 10659
rect 13737 10625 13771 10659
rect 13829 10625 13863 10659
rect 14105 10625 14139 10659
rect 18245 10625 18279 10659
rect 2237 10557 2271 10591
rect 14289 10557 14323 10591
rect 1501 10421 1535 10455
rect 4997 10421 5031 10455
rect 18429 10421 18463 10455
rect 17601 10217 17635 10251
rect 17785 10217 17819 10251
rect 5089 10149 5123 10183
rect 15025 10149 15059 10183
rect 1685 10081 1719 10115
rect 10701 10081 10735 10115
rect 11805 10081 11839 10115
rect 17417 10081 17451 10115
rect 17877 10081 17911 10115
rect 1501 10013 1535 10047
rect 1869 10013 1903 10047
rect 2053 10013 2087 10047
rect 4905 10013 4939 10047
rect 10609 10013 10643 10047
rect 11437 10013 11471 10047
rect 11713 10013 11747 10047
rect 14657 10013 14691 10047
rect 15117 10013 15151 10047
rect 16589 10013 16623 10047
rect 16957 10013 16991 10047
rect 17785 10013 17819 10047
rect 18245 10013 18279 10047
rect 14749 9945 14783 9979
rect 15393 9945 15427 9979
rect 16405 9945 16439 9979
rect 1961 9877 1995 9911
rect 10977 9877 11011 9911
rect 14473 9877 14507 9911
rect 14841 9877 14875 9911
rect 1593 9673 1627 9707
rect 5381 9673 5415 9707
rect 3249 9605 3283 9639
rect 5181 9605 5215 9639
rect 18429 9605 18463 9639
rect 1409 9537 1443 9571
rect 2053 9537 2087 9571
rect 2329 9537 2363 9571
rect 2421 9537 2455 9571
rect 2973 9537 3007 9571
rect 3157 9537 3191 9571
rect 3341 9537 3375 9571
rect 6009 9537 6043 9571
rect 16209 9535 16243 9569
rect 16681 9537 16715 9571
rect 16865 9537 16899 9571
rect 17969 9537 18003 9571
rect 18337 9537 18371 9571
rect 5733 9469 5767 9503
rect 5825 9469 5859 9503
rect 5917 9469 5951 9503
rect 16037 9469 16071 9503
rect 18245 9469 18279 9503
rect 3525 9401 3559 9435
rect 5549 9401 5583 9435
rect 18061 9401 18095 9435
rect 2145 9333 2179 9367
rect 2605 9333 2639 9367
rect 5365 9333 5399 9367
rect 6193 9333 6227 9367
rect 16405 9333 16439 9367
rect 16773 9333 16807 9367
rect 2145 9129 2179 9163
rect 17693 9129 17727 9163
rect 17785 9129 17819 9163
rect 17969 9061 18003 9095
rect 17877 8993 17911 9027
rect 1961 8925 1995 8959
rect 2145 8925 2179 8959
rect 8953 8925 8987 8959
rect 9149 8925 9183 8959
rect 14749 8925 14783 8959
rect 15025 8925 15059 8959
rect 17601 8925 17635 8959
rect 17969 8925 18003 8959
rect 18153 8925 18187 8959
rect 18245 8925 18279 8959
rect 9045 8789 9079 8823
rect 14381 8789 14415 8823
rect 18429 8789 18463 8823
rect 4169 8585 4203 8619
rect 7113 8585 7147 8619
rect 12449 8585 12483 8619
rect 14197 8585 14231 8619
rect 14565 8585 14599 8619
rect 6653 8517 6687 8551
rect 16405 8517 16439 8551
rect 3617 8449 3651 8483
rect 3709 8449 3743 8483
rect 3893 8449 3927 8483
rect 3985 8449 4019 8483
rect 4537 8449 4571 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 6929 8449 6963 8483
rect 7021 8449 7055 8483
rect 7573 8449 7607 8483
rect 10149 8449 10183 8483
rect 12357 8449 12391 8483
rect 12541 8449 12575 8483
rect 14105 8449 14139 8483
rect 14381 8449 14415 8483
rect 16129 8449 16163 8483
rect 16221 8449 16255 8483
rect 1409 8381 1443 8415
rect 1685 8381 1719 8415
rect 4445 8381 4479 8415
rect 7205 8381 7239 8415
rect 7297 8381 7331 8415
rect 3433 8313 3467 8347
rect 9689 8313 9723 8347
rect 4445 8245 4479 8279
rect 6377 8245 6411 8279
rect 7481 8245 7515 8279
rect 9873 8245 9907 8279
rect 16129 8245 16163 8279
rect 2513 8041 2547 8075
rect 3249 8041 3283 8075
rect 17877 8041 17911 8075
rect 2697 7905 2731 7939
rect 8125 7905 8159 7939
rect 2053 7837 2087 7871
rect 2329 7837 2363 7871
rect 2605 7837 2639 7871
rect 2789 7837 2823 7871
rect 3433 7837 3467 7871
rect 3985 7837 4019 7871
rect 4353 7837 4387 7871
rect 4721 7837 4755 7871
rect 8033 7837 8067 7871
rect 8309 7837 8343 7871
rect 8401 7837 8435 7871
rect 17693 7837 17727 7871
rect 3617 7769 3651 7803
rect 4905 7769 4939 7803
rect 2145 7701 2179 7735
rect 8585 7701 8619 7735
rect 13353 7497 13387 7531
rect 14381 7497 14415 7531
rect 1685 7429 1719 7463
rect 8125 7429 8159 7463
rect 13553 7429 13587 7463
rect 1501 7361 1535 7395
rect 7941 7361 7975 7395
rect 8033 7361 8067 7395
rect 8309 7361 8343 7395
rect 8401 7361 8435 7395
rect 13829 7361 13863 7395
rect 14105 7361 14139 7395
rect 14197 7361 14231 7395
rect 13921 7293 13955 7327
rect 16313 7293 16347 7327
rect 15945 7225 15979 7259
rect 7757 7157 7791 7191
rect 13185 7157 13219 7191
rect 13369 7157 13403 7191
rect 15853 7157 15887 7191
rect 9413 6953 9447 6987
rect 2605 6817 2639 6851
rect 5089 6817 5123 6851
rect 16221 6817 16255 6851
rect 2789 6749 2823 6783
rect 4997 6749 5031 6783
rect 5181 6749 5215 6783
rect 9689 6749 9723 6783
rect 9965 6749 9999 6783
rect 10057 6749 10091 6783
rect 12449 6749 12483 6783
rect 12541 6749 12575 6783
rect 12633 6749 12667 6783
rect 15301 6749 15335 6783
rect 15761 6749 15795 6783
rect 16037 6749 16071 6783
rect 16773 6749 16807 6783
rect 18245 6749 18279 6783
rect 2973 6681 3007 6715
rect 3157 6681 3191 6715
rect 9597 6681 9631 6715
rect 9873 6681 9907 6715
rect 2881 6613 2915 6647
rect 9229 6613 9263 6647
rect 9397 6613 9431 6647
rect 10241 6613 10275 6647
rect 18429 6613 18463 6647
rect 2053 6409 2087 6443
rect 6644 6409 6678 6443
rect 10425 6409 10459 6443
rect 18245 6409 18279 6443
rect 1409 6341 1443 6375
rect 1625 6341 1659 6375
rect 13737 6341 13771 6375
rect 1869 6273 1903 6307
rect 6377 6273 6411 6307
rect 7021 6273 7055 6307
rect 9965 6273 9999 6307
rect 16221 6273 16255 6307
rect 18521 6273 18555 6307
rect 13277 6205 13311 6239
rect 16129 6205 16163 6239
rect 18245 6205 18279 6239
rect 1777 6137 1811 6171
rect 13369 6137 13403 6171
rect 15853 6137 15887 6171
rect 18429 6137 18463 6171
rect 1593 6069 1627 6103
rect 6653 6069 6687 6103
rect 10241 6069 10275 6103
rect 4261 5865 4295 5899
rect 4445 5865 4479 5899
rect 14749 5865 14783 5899
rect 16773 5865 16807 5899
rect 11529 5729 11563 5763
rect 14105 5729 14139 5763
rect 11897 5661 11931 5695
rect 12173 5661 12207 5695
rect 12909 5661 12943 5695
rect 13461 5661 13495 5695
rect 14197 5661 14231 5695
rect 14381 5661 14415 5695
rect 14657 5661 14691 5695
rect 14841 5661 14875 5695
rect 16129 5661 16163 5695
rect 16405 5661 16439 5695
rect 16865 5661 16899 5695
rect 4077 5593 4111 5627
rect 4293 5593 4327 5627
rect 16589 5593 16623 5627
rect 13185 5525 13219 5559
rect 14565 5525 14599 5559
rect 16221 5525 16255 5559
rect 1593 5321 1627 5355
rect 2513 5321 2547 5355
rect 5273 5321 5307 5355
rect 8033 5321 8067 5355
rect 15393 5321 15427 5355
rect 7849 5253 7883 5287
rect 11989 5253 12023 5287
rect 13001 5253 13035 5287
rect 1409 5185 1443 5219
rect 2237 5185 2271 5219
rect 7757 5185 7791 5219
rect 8125 5185 8159 5219
rect 12633 5185 12667 5219
rect 12817 5185 12851 5219
rect 13369 5185 13403 5219
rect 13461 5185 13495 5219
rect 13737 5185 13771 5219
rect 15209 5185 15243 5219
rect 15393 5185 15427 5219
rect 4813 5117 4847 5151
rect 7941 5117 7975 5151
rect 13185 5117 13219 5151
rect 5181 5049 5215 5083
rect 12081 4981 12115 5015
rect 13645 4981 13679 5015
rect 14105 4777 14139 4811
rect 14289 4777 14323 4811
rect 16681 4777 16715 4811
rect 16773 4777 16807 4811
rect 10057 4709 10091 4743
rect 12081 4709 12115 4743
rect 12449 4709 12483 4743
rect 9229 4641 9263 4675
rect 9321 4641 9355 4675
rect 9413 4641 9447 4675
rect 12541 4641 12575 4675
rect 9137 4573 9171 4607
rect 10885 4573 10919 4607
rect 11069 4573 11103 4607
rect 12265 4573 12299 4607
rect 14657 4573 14691 4607
rect 15669 4573 15703 4607
rect 16037 4573 16071 4607
rect 16129 4573 16163 4607
rect 16497 4573 16531 4607
rect 16773 4573 16807 4607
rect 16957 4573 16991 4607
rect 16313 4505 16347 4539
rect 16405 4505 16439 4539
rect 8953 4437 8987 4471
rect 14289 4437 14323 4471
rect 10057 4233 10091 4267
rect 10149 4233 10183 4267
rect 3157 4165 3191 4199
rect 10241 4165 10275 4199
rect 14533 4165 14567 4199
rect 14749 4165 14783 4199
rect 17509 4165 17543 4199
rect 1409 4097 1443 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 17325 4097 17359 4131
rect 18245 4097 18279 4131
rect 17693 4029 17727 4063
rect 1593 3961 1627 3995
rect 5825 3961 5859 3995
rect 9873 3961 9907 3995
rect 3065 3893 3099 3927
rect 10425 3893 10459 3927
rect 14381 3893 14415 3927
rect 14565 3893 14599 3927
rect 18429 3893 18463 3927
rect 3893 3689 3927 3723
rect 4353 3689 4387 3723
rect 15301 3689 15335 3723
rect 9137 3621 9171 3655
rect 14657 3553 14691 3587
rect 3801 3485 3835 3519
rect 4077 3485 4111 3519
rect 9321 3485 9355 3519
rect 9413 3485 9447 3519
rect 15025 3485 15059 3519
rect 15117 3485 15151 3519
rect 9137 3417 9171 3451
rect 1685 3077 1719 3111
rect 4077 3077 4111 3111
rect 12265 3077 12299 3111
rect 12357 3077 12391 3111
rect 14289 3077 14323 3111
rect 14473 3077 14507 3111
rect 1501 3009 1535 3043
rect 1869 3009 1903 3043
rect 2145 3009 2179 3043
rect 2329 3009 2363 3043
rect 3801 3009 3835 3043
rect 3893 3009 3927 3043
rect 8953 3009 8987 3043
rect 9137 3009 9171 3043
rect 9229 3009 9263 3043
rect 10977 3009 11011 3043
rect 11161 3009 11195 3043
rect 11989 3009 12023 3043
rect 12137 3009 12171 3043
rect 12495 3009 12529 3043
rect 14565 3009 14599 3043
rect 11345 2941 11379 2975
rect 2053 2873 2087 2907
rect 14289 2873 14323 2907
rect 2329 2805 2363 2839
rect 4077 2805 4111 2839
rect 12633 2805 12667 2839
rect 4169 2601 4203 2635
rect 9045 2601 9079 2635
rect 17877 2601 17911 2635
rect 1869 2533 1903 2567
rect 10425 2533 10459 2567
rect 17693 2533 17727 2567
rect 16957 2465 16991 2499
rect 1685 2397 1719 2431
rect 1777 2397 1811 2431
rect 2329 2397 2363 2431
rect 8953 2397 8987 2431
rect 9137 2397 9171 2431
rect 15761 2397 15795 2431
rect 16773 2397 16807 2431
rect 18245 2397 18279 2431
rect 3893 2329 3927 2363
rect 10149 2329 10183 2363
rect 15945 2329 15979 2363
rect 16129 2329 16163 2363
rect 17845 2329 17879 2363
rect 18061 2329 18095 2363
rect 18429 2261 18463 2295
<< metal1 >>
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 18138 17660 18144 17672
rect 5500 17632 18144 17660
rect 5500 17620 5506 17632
rect 18138 17620 18144 17632
rect 18196 17620 18202 17672
rect 13262 17552 13268 17604
rect 13320 17592 13326 17604
rect 16574 17592 16580 17604
rect 13320 17564 16580 17592
rect 13320 17552 13326 17564
rect 16574 17552 16580 17564
rect 16632 17552 16638 17604
rect 9306 17484 9312 17536
rect 9364 17524 9370 17536
rect 18230 17524 18236 17536
rect 9364 17496 18236 17524
rect 9364 17484 9370 17496
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 1104 17434 18860 17456
rect 1104 17382 2610 17434
rect 2662 17382 2674 17434
rect 2726 17382 2738 17434
rect 2790 17382 2802 17434
rect 2854 17382 2866 17434
rect 2918 17382 7610 17434
rect 7662 17382 7674 17434
rect 7726 17382 7738 17434
rect 7790 17382 7802 17434
rect 7854 17382 7866 17434
rect 7918 17382 12610 17434
rect 12662 17382 12674 17434
rect 12726 17382 12738 17434
rect 12790 17382 12802 17434
rect 12854 17382 12866 17434
rect 12918 17382 17610 17434
rect 17662 17382 17674 17434
rect 17726 17382 17738 17434
rect 17790 17382 17802 17434
rect 17854 17382 17866 17434
rect 17918 17382 18860 17434
rect 1104 17360 18860 17382
rect 13262 17320 13268 17332
rect 2884 17292 13268 17320
rect 1854 17212 1860 17264
rect 1912 17212 1918 17264
rect 2884 17261 2912 17292
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 17954 17280 17960 17332
rect 18012 17320 18018 17332
rect 18417 17323 18475 17329
rect 18417 17320 18429 17323
rect 18012 17292 18429 17320
rect 18012 17280 18018 17292
rect 18417 17289 18429 17292
rect 18463 17289 18475 17323
rect 18417 17283 18475 17289
rect 2869 17255 2927 17261
rect 2869 17221 2881 17255
rect 2915 17221 2927 17255
rect 10502 17252 10508 17264
rect 2869 17215 2927 17221
rect 5276 17224 10508 17252
rect 842 17144 848 17196
rect 900 17184 906 17196
rect 1489 17187 1547 17193
rect 1489 17184 1501 17187
rect 900 17156 1501 17184
rect 900 17144 906 17156
rect 1489 17153 1501 17156
rect 1535 17153 1547 17187
rect 1489 17147 1547 17153
rect 2498 17144 2504 17196
rect 2556 17144 2562 17196
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 5074 17184 5080 17196
rect 2823 17156 5080 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 5074 17144 5080 17156
rect 5132 17184 5138 17196
rect 5276 17184 5304 17224
rect 10502 17212 10508 17224
rect 10560 17252 10566 17264
rect 13630 17252 13636 17264
rect 10560 17224 13636 17252
rect 10560 17212 10566 17224
rect 13630 17212 13636 17224
rect 13688 17212 13694 17264
rect 13722 17212 13728 17264
rect 13780 17252 13786 17264
rect 13780 17224 15332 17252
rect 13780 17212 13786 17224
rect 5132 17156 5304 17184
rect 5353 17187 5411 17193
rect 5132 17144 5138 17156
rect 5353 17153 5365 17187
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 5368 17116 5396 17147
rect 8846 17144 8852 17196
rect 8904 17184 8910 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 8904 17156 14749 17184
rect 8904 17144 8910 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 2746 17088 5396 17116
rect 1673 17051 1731 17057
rect 1673 17017 1685 17051
rect 1719 17048 1731 17051
rect 2314 17048 2320 17060
rect 1719 17020 2320 17048
rect 1719 17017 1731 17020
rect 1673 17011 1731 17017
rect 2314 17008 2320 17020
rect 2372 17008 2378 17060
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 1949 16983 2007 16989
rect 1949 16980 1961 16983
rect 1452 16952 1961 16980
rect 1452 16940 1458 16952
rect 1949 16949 1961 16952
rect 1995 16980 2007 16983
rect 2746 16980 2774 17088
rect 10042 17076 10048 17128
rect 10100 17116 10106 17128
rect 14458 17116 14464 17128
rect 10100 17088 14464 17116
rect 10100 17076 10106 17088
rect 14458 17076 14464 17088
rect 14516 17076 14522 17128
rect 15194 17076 15200 17128
rect 15252 17076 15258 17128
rect 15304 17116 15332 17224
rect 15565 17187 15623 17193
rect 15565 17153 15577 17187
rect 15611 17184 15623 17187
rect 16390 17184 16396 17196
rect 15611 17156 16396 17184
rect 15611 17153 15623 17156
rect 15565 17147 15623 17153
rect 16390 17144 16396 17156
rect 16448 17144 16454 17196
rect 18230 17144 18236 17196
rect 18288 17144 18294 17196
rect 16025 17119 16083 17125
rect 16025 17116 16037 17119
rect 15304 17088 16037 17116
rect 16025 17085 16037 17088
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 4154 17008 4160 17060
rect 4212 17048 4218 17060
rect 10226 17048 10232 17060
rect 4212 17020 10232 17048
rect 4212 17008 4218 17020
rect 10226 17008 10232 17020
rect 10284 17008 10290 17060
rect 11790 17008 11796 17060
rect 11848 17048 11854 17060
rect 15654 17048 15660 17060
rect 11848 17020 15660 17048
rect 11848 17008 11854 17020
rect 15654 17008 15660 17020
rect 15712 17008 15718 17060
rect 1995 16952 2774 16980
rect 1995 16949 2007 16952
rect 1949 16943 2007 16949
rect 5258 16940 5264 16992
rect 5316 16940 5322 16992
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 9766 16980 9772 16992
rect 5592 16952 9772 16980
rect 5592 16940 5598 16952
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10778 16940 10784 16992
rect 10836 16980 10842 16992
rect 14642 16980 14648 16992
rect 10836 16952 14648 16980
rect 10836 16940 10842 16952
rect 14642 16940 14648 16952
rect 14700 16940 14706 16992
rect 1104 16890 18860 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 6950 16890
rect 7002 16838 7014 16890
rect 7066 16838 7078 16890
rect 7130 16838 7142 16890
rect 7194 16838 7206 16890
rect 7258 16838 11950 16890
rect 12002 16838 12014 16890
rect 12066 16838 12078 16890
rect 12130 16838 12142 16890
rect 12194 16838 12206 16890
rect 12258 16838 16950 16890
rect 17002 16838 17014 16890
rect 17066 16838 17078 16890
rect 17130 16838 17142 16890
rect 17194 16838 17206 16890
rect 17258 16838 18860 16890
rect 1104 16816 18860 16838
rect 4982 16736 4988 16788
rect 5040 16776 5046 16788
rect 5442 16776 5448 16788
rect 5040 16748 5448 16776
rect 5040 16736 5046 16748
rect 5442 16736 5448 16748
rect 5500 16776 5506 16788
rect 5537 16779 5595 16785
rect 5537 16776 5549 16779
rect 5500 16748 5549 16776
rect 5500 16736 5506 16748
rect 5537 16745 5549 16748
rect 5583 16745 5595 16779
rect 8294 16776 8300 16788
rect 5537 16739 5595 16745
rect 5736 16748 8300 16776
rect 4154 16668 4160 16720
rect 4212 16668 4218 16720
rect 5534 16532 5540 16584
rect 5592 16532 5598 16584
rect 5736 16581 5764 16748
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 9490 16736 9496 16788
rect 9548 16776 9554 16788
rect 9858 16776 9864 16788
rect 9548 16748 9864 16776
rect 9548 16736 9554 16748
rect 9858 16736 9864 16748
rect 9916 16776 9922 16788
rect 11238 16776 11244 16788
rect 9916 16748 9996 16776
rect 9916 16736 9922 16748
rect 6546 16668 6552 16720
rect 6604 16708 6610 16720
rect 9674 16708 9680 16720
rect 6604 16680 9680 16708
rect 6604 16668 6610 16680
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 5721 16575 5779 16581
rect 5721 16541 5733 16575
rect 5767 16541 5779 16575
rect 5721 16535 5779 16541
rect 3694 16464 3700 16516
rect 3752 16504 3758 16516
rect 3789 16507 3847 16513
rect 3789 16504 3801 16507
rect 3752 16476 3801 16504
rect 3752 16464 3758 16476
rect 3789 16473 3801 16476
rect 3835 16473 3847 16507
rect 3789 16467 3847 16473
rect 4249 16439 4307 16445
rect 4249 16405 4261 16439
rect 4295 16436 4307 16439
rect 6656 16436 6684 16603
rect 6822 16600 6828 16652
rect 6880 16600 6886 16652
rect 6932 16649 6960 16680
rect 9674 16668 9680 16680
rect 9732 16668 9738 16720
rect 9968 16717 9996 16748
rect 10520 16748 11244 16776
rect 9953 16711 10011 16717
rect 9953 16677 9965 16711
rect 9999 16677 10011 16711
rect 9953 16671 10011 16677
rect 6917 16643 6975 16649
rect 6917 16609 6929 16643
rect 6963 16609 6975 16643
rect 10520 16640 10548 16748
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 15654 16736 15660 16788
rect 15712 16736 15718 16788
rect 18141 16779 18199 16785
rect 16224 16748 18092 16776
rect 10597 16711 10655 16717
rect 10597 16677 10609 16711
rect 10643 16677 10655 16711
rect 10597 16671 10655 16677
rect 6917 16603 6975 16609
rect 8496 16612 10548 16640
rect 8392 16584 8444 16590
rect 6730 16532 6736 16584
rect 6788 16532 6794 16584
rect 8496 16581 8524 16612
rect 8481 16575 8539 16581
rect 8481 16541 8493 16575
rect 8527 16541 8539 16575
rect 8481 16535 8539 16541
rect 8754 16532 8760 16584
rect 8812 16572 8818 16584
rect 8941 16575 8999 16581
rect 8941 16572 8953 16575
rect 8812 16544 8953 16572
rect 8812 16532 8818 16544
rect 8941 16541 8953 16544
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 9122 16532 9128 16584
rect 9180 16532 9186 16584
rect 9582 16532 9588 16584
rect 9640 16572 9646 16584
rect 9677 16575 9735 16581
rect 9677 16572 9689 16575
rect 9640 16544 9689 16572
rect 9640 16532 9646 16544
rect 9677 16541 9689 16544
rect 9723 16572 9735 16575
rect 10042 16572 10048 16584
rect 9723 16544 10048 16572
rect 9723 16541 9735 16544
rect 9677 16535 9735 16541
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 10318 16532 10324 16584
rect 10376 16532 10382 16584
rect 10612 16572 10640 16671
rect 13906 16668 13912 16720
rect 13964 16708 13970 16720
rect 14921 16711 14979 16717
rect 13964 16680 14780 16708
rect 13964 16668 13970 16680
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 13541 16643 13599 16649
rect 13541 16640 13553 16643
rect 10744 16612 13553 16640
rect 10744 16600 10750 16612
rect 13541 16609 13553 16612
rect 13587 16609 13599 16643
rect 13541 16603 13599 16609
rect 13630 16600 13636 16652
rect 13688 16640 13694 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13688 16612 14105 16640
rect 13688 16600 13694 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 14274 16600 14280 16652
rect 14332 16640 14338 16652
rect 14332 16612 14596 16640
rect 14332 16600 14338 16612
rect 10870 16572 10876 16584
rect 10612 16544 10876 16572
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 12805 16575 12863 16581
rect 12805 16541 12817 16575
rect 12851 16541 12863 16575
rect 12805 16535 12863 16541
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16541 13139 16575
rect 13081 16535 13139 16541
rect 8392 16526 8444 16532
rect 7374 16464 7380 16516
rect 7432 16504 7438 16516
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 7432 16476 7481 16504
rect 7432 16464 7438 16476
rect 7469 16473 7481 16476
rect 7515 16473 7527 16507
rect 7469 16467 7527 16473
rect 9950 16464 9956 16516
rect 10008 16464 10014 16516
rect 10594 16464 10600 16516
rect 10652 16464 10658 16516
rect 12434 16464 12440 16516
rect 12492 16504 12498 16516
rect 12820 16504 12848 16535
rect 12492 16476 12848 16504
rect 13096 16504 13124 16535
rect 14458 16532 14464 16584
rect 14516 16532 14522 16584
rect 14568 16572 14596 16612
rect 14642 16600 14648 16652
rect 14700 16600 14706 16652
rect 14752 16640 14780 16680
rect 14921 16677 14933 16711
rect 14967 16708 14979 16711
rect 16224 16708 16252 16748
rect 16758 16708 16764 16720
rect 14967 16680 16252 16708
rect 16316 16680 16764 16708
rect 14967 16677 14979 16680
rect 14921 16671 14979 16677
rect 15749 16643 15807 16649
rect 14752 16612 14964 16640
rect 14936 16581 14964 16612
rect 15749 16609 15761 16643
rect 15795 16640 15807 16643
rect 16316 16640 16344 16680
rect 16758 16668 16764 16680
rect 16816 16668 16822 16720
rect 18064 16708 18092 16748
rect 18141 16745 18153 16779
rect 18187 16776 18199 16779
rect 18322 16776 18328 16788
rect 18187 16748 18328 16776
rect 18187 16745 18199 16748
rect 18141 16739 18199 16745
rect 18322 16736 18328 16748
rect 18380 16736 18386 16788
rect 18506 16708 18512 16720
rect 18064 16680 18512 16708
rect 18506 16668 18512 16680
rect 18564 16668 18570 16720
rect 17037 16643 17095 16649
rect 15795 16612 16344 16640
rect 16408 16612 16804 16640
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 14737 16575 14795 16581
rect 14737 16572 14749 16575
rect 14568 16544 14749 16572
rect 14737 16541 14749 16544
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 14921 16575 14979 16581
rect 14921 16541 14933 16575
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 15010 16532 15016 16584
rect 15068 16532 15074 16584
rect 15194 16532 15200 16584
rect 15252 16532 15258 16584
rect 15657 16575 15715 16581
rect 15657 16572 15669 16575
rect 15304 16544 15669 16572
rect 13262 16504 13268 16516
rect 13096 16476 13268 16504
rect 12492 16464 12498 16476
rect 13262 16464 13268 16476
rect 13320 16464 13326 16516
rect 14182 16464 14188 16516
rect 14240 16464 14246 16516
rect 15105 16507 15163 16513
rect 15105 16504 15117 16507
rect 14292 16476 15117 16504
rect 4295 16408 6684 16436
rect 7101 16439 7159 16445
rect 4295 16405 4307 16408
rect 4249 16399 4307 16405
rect 7101 16405 7113 16439
rect 7147 16436 7159 16439
rect 7282 16436 7288 16448
rect 7147 16408 7288 16436
rect 7147 16405 7159 16408
rect 7101 16399 7159 16405
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 9030 16396 9036 16448
rect 9088 16396 9094 16448
rect 9769 16439 9827 16445
rect 9769 16405 9781 16439
rect 9815 16436 9827 16439
rect 10134 16436 10140 16448
rect 9815 16408 10140 16436
rect 9815 16405 9827 16408
rect 9769 16399 9827 16405
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 10318 16396 10324 16448
rect 10376 16436 10382 16448
rect 10413 16439 10471 16445
rect 10413 16436 10425 16439
rect 10376 16408 10425 16436
rect 10376 16396 10382 16408
rect 10413 16405 10425 16408
rect 10459 16405 10471 16439
rect 10413 16399 10471 16405
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 14292 16436 14320 16476
rect 15105 16473 15117 16476
rect 15151 16473 15163 16507
rect 15105 16467 15163 16473
rect 11204 16408 14320 16436
rect 11204 16396 11210 16408
rect 14918 16396 14924 16448
rect 14976 16436 14982 16448
rect 15304 16436 15332 16544
rect 15657 16541 15669 16544
rect 15703 16541 15715 16575
rect 15657 16535 15715 16541
rect 15378 16464 15384 16516
rect 15436 16504 15442 16516
rect 16408 16504 16436 16612
rect 16485 16575 16543 16581
rect 16485 16541 16497 16575
rect 16531 16541 16543 16575
rect 16485 16535 16543 16541
rect 16577 16575 16635 16581
rect 16577 16541 16589 16575
rect 16623 16572 16635 16575
rect 16666 16572 16672 16584
rect 16623 16544 16672 16572
rect 16623 16541 16635 16544
rect 16577 16535 16635 16541
rect 15436 16476 16436 16504
rect 16500 16504 16528 16535
rect 16666 16532 16672 16544
rect 16724 16532 16730 16584
rect 16776 16581 16804 16612
rect 17037 16609 17049 16643
rect 17083 16640 17095 16643
rect 18782 16640 18788 16652
rect 17083 16612 18788 16640
rect 17083 16609 17095 16612
rect 17037 16603 17095 16609
rect 18782 16600 18788 16612
rect 18840 16600 18846 16652
rect 16761 16575 16819 16581
rect 16761 16541 16773 16575
rect 16807 16541 16819 16575
rect 16761 16535 16819 16541
rect 16850 16532 16856 16584
rect 16908 16532 16914 16584
rect 16942 16532 16948 16584
rect 17000 16572 17006 16584
rect 17589 16575 17647 16581
rect 17589 16572 17601 16575
rect 17000 16544 17601 16572
rect 17000 16532 17006 16544
rect 17589 16541 17601 16544
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 17310 16504 17316 16516
rect 16500 16476 17316 16504
rect 15436 16464 15442 16476
rect 17310 16464 17316 16476
rect 17368 16464 17374 16516
rect 17402 16464 17408 16516
rect 17460 16504 17466 16516
rect 18325 16507 18383 16513
rect 18325 16504 18337 16507
rect 17460 16476 18337 16504
rect 17460 16464 17466 16476
rect 18325 16473 18337 16476
rect 18371 16473 18383 16507
rect 18325 16467 18383 16473
rect 14976 16408 15332 16436
rect 14976 16396 14982 16408
rect 15930 16396 15936 16448
rect 15988 16436 15994 16448
rect 16025 16439 16083 16445
rect 16025 16436 16037 16439
rect 15988 16408 16037 16436
rect 15988 16396 15994 16408
rect 16025 16405 16037 16408
rect 16071 16405 16083 16439
rect 16025 16399 16083 16405
rect 17494 16396 17500 16448
rect 17552 16436 17558 16448
rect 17773 16439 17831 16445
rect 17773 16436 17785 16439
rect 17552 16408 17785 16436
rect 17552 16396 17558 16408
rect 17773 16405 17785 16408
rect 17819 16405 17831 16439
rect 17773 16399 17831 16405
rect 17954 16396 17960 16448
rect 18012 16396 18018 16448
rect 18125 16439 18183 16445
rect 18125 16405 18137 16439
rect 18171 16436 18183 16439
rect 18414 16436 18420 16448
rect 18171 16408 18420 16436
rect 18171 16405 18183 16408
rect 18125 16399 18183 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 1104 16346 18860 16368
rect 1104 16294 2610 16346
rect 2662 16294 2674 16346
rect 2726 16294 2738 16346
rect 2790 16294 2802 16346
rect 2854 16294 2866 16346
rect 2918 16294 7610 16346
rect 7662 16294 7674 16346
rect 7726 16294 7738 16346
rect 7790 16294 7802 16346
rect 7854 16294 7866 16346
rect 7918 16294 12610 16346
rect 12662 16294 12674 16346
rect 12726 16294 12738 16346
rect 12790 16294 12802 16346
rect 12854 16294 12866 16346
rect 12918 16294 17610 16346
rect 17662 16294 17674 16346
rect 17726 16294 17738 16346
rect 17790 16294 17802 16346
rect 17854 16294 17866 16346
rect 17918 16294 18860 16346
rect 1104 16272 18860 16294
rect 1673 16235 1731 16241
rect 1673 16201 1685 16235
rect 1719 16232 1731 16235
rect 2958 16232 2964 16244
rect 1719 16204 2964 16232
rect 1719 16201 1731 16204
rect 1673 16195 1731 16201
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 5626 16192 5632 16244
rect 5684 16232 5690 16244
rect 9490 16232 9496 16244
rect 5684 16204 9496 16232
rect 5684 16192 5690 16204
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 13170 16232 13176 16244
rect 11572 16204 13176 16232
rect 11572 16192 11578 16204
rect 13170 16192 13176 16204
rect 13228 16192 13234 16244
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 17865 16235 17923 16241
rect 17865 16232 17877 16235
rect 15528 16204 17877 16232
rect 15528 16192 15534 16204
rect 17865 16201 17877 16204
rect 17911 16201 17923 16235
rect 17865 16195 17923 16201
rect 1026 16124 1032 16176
rect 1084 16164 1090 16176
rect 1949 16167 2007 16173
rect 1949 16164 1961 16167
rect 1084 16136 1961 16164
rect 1084 16124 1090 16136
rect 1949 16133 1961 16136
rect 1995 16133 2007 16167
rect 4062 16164 4068 16176
rect 1949 16127 2007 16133
rect 2746 16136 4068 16164
rect 1489 16099 1547 16105
rect 1489 16065 1501 16099
rect 1535 16096 1547 16099
rect 1578 16096 1584 16108
rect 1535 16068 1584 16096
rect 1535 16065 1547 16068
rect 1489 16059 1547 16065
rect 1578 16056 1584 16068
rect 1636 16056 1642 16108
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 2498 16096 2504 16108
rect 1811 16068 2504 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 2498 16056 2504 16068
rect 2556 16096 2562 16108
rect 2746 16096 2774 16136
rect 4062 16124 4068 16136
rect 4120 16164 4126 16176
rect 9398 16164 9404 16176
rect 4120 16136 9404 16164
rect 4120 16124 4126 16136
rect 9398 16124 9404 16136
rect 9456 16124 9462 16176
rect 9858 16124 9864 16176
rect 9916 16164 9922 16176
rect 9916 16136 11928 16164
rect 9916 16124 9922 16136
rect 2556 16068 2774 16096
rect 2556 16056 2562 16068
rect 3050 16056 3056 16108
rect 3108 16056 3114 16108
rect 3142 16056 3148 16108
rect 3200 16096 3206 16108
rect 3513 16099 3571 16105
rect 3513 16096 3525 16099
rect 3200 16068 3525 16096
rect 3200 16056 3206 16068
rect 3513 16065 3525 16068
rect 3559 16065 3571 16099
rect 3513 16059 3571 16065
rect 9585 16099 9643 16105
rect 9585 16065 9597 16099
rect 9631 16096 9643 16099
rect 9950 16096 9956 16108
rect 9631 16068 9956 16096
rect 9631 16065 9643 16068
rect 9585 16059 9643 16065
rect 9950 16056 9956 16068
rect 10008 16056 10014 16108
rect 10042 16056 10048 16108
rect 10100 16096 10106 16108
rect 11900 16105 11928 16136
rect 11974 16124 11980 16176
rect 12032 16164 12038 16176
rect 12805 16167 12863 16173
rect 12805 16164 12817 16167
rect 12032 16136 12817 16164
rect 12032 16124 12038 16136
rect 12805 16133 12817 16136
rect 12851 16164 12863 16167
rect 18874 16164 18880 16176
rect 12851 16136 18880 16164
rect 12851 16133 12863 16136
rect 12805 16127 12863 16133
rect 18874 16124 18880 16136
rect 18932 16124 18938 16176
rect 11793 16099 11851 16105
rect 11793 16096 11805 16099
rect 10100 16068 11805 16096
rect 10100 16056 10106 16068
rect 11793 16065 11805 16068
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 12986 16056 12992 16108
rect 13044 16096 13050 16108
rect 13173 16099 13231 16105
rect 13173 16096 13185 16099
rect 13044 16068 13185 16096
rect 13044 16056 13050 16068
rect 13173 16065 13185 16068
rect 13219 16065 13231 16099
rect 13173 16059 13231 16065
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 13320 16068 13369 16096
rect 13320 16056 13326 16068
rect 13357 16065 13369 16068
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 13446 16056 13452 16108
rect 13504 16096 13510 16108
rect 13541 16099 13599 16105
rect 13541 16096 13553 16099
rect 13504 16068 13553 16096
rect 13504 16056 13510 16068
rect 13541 16065 13553 16068
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 14550 16056 14556 16108
rect 14608 16096 14614 16108
rect 17773 16099 17831 16105
rect 17773 16096 17785 16099
rect 14608 16068 17785 16096
rect 14608 16056 14614 16068
rect 17773 16065 17785 16068
rect 17819 16065 17831 16099
rect 17773 16059 17831 16065
rect 18138 16056 18144 16108
rect 18196 16096 18202 16108
rect 18233 16099 18291 16105
rect 18233 16096 18245 16099
rect 18196 16068 18245 16096
rect 18196 16056 18202 16068
rect 18233 16065 18245 16068
rect 18279 16096 18291 16099
rect 18598 16096 18604 16108
rect 18279 16068 18604 16096
rect 18279 16065 18291 16068
rect 18233 16059 18291 16065
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 4341 16031 4399 16037
rect 4341 15997 4353 16031
rect 4387 16028 4399 16031
rect 4798 16028 4804 16040
rect 4387 16000 4804 16028
rect 4387 15997 4399 16000
rect 4341 15991 4399 15997
rect 4798 15988 4804 16000
rect 4856 15988 4862 16040
rect 9398 15988 9404 16040
rect 9456 15988 9462 16040
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 1486 15920 1492 15972
rect 1544 15920 1550 15972
rect 2133 15963 2191 15969
rect 2133 15929 2145 15963
rect 2179 15960 2191 15963
rect 9214 15960 9220 15972
rect 2179 15932 9220 15960
rect 2179 15929 2191 15932
rect 2133 15923 2191 15929
rect 9214 15920 9220 15932
rect 9272 15920 9278 15972
rect 9508 15960 9536 15991
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 10962 16028 10968 16040
rect 9732 16000 10968 16028
rect 9732 15988 9738 16000
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 11330 15988 11336 16040
rect 11388 16028 11394 16040
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 11388 16000 12081 16028
rect 11388 15988 11394 16000
rect 12069 15997 12081 16000
rect 12115 15997 12127 16031
rect 12069 15991 12127 15997
rect 12894 15988 12900 16040
rect 12952 16028 12958 16040
rect 14918 16028 14924 16040
rect 12952 16000 14924 16028
rect 12952 15988 12958 16000
rect 14918 15988 14924 16000
rect 14976 15988 14982 16040
rect 11348 15960 11376 15988
rect 9508 15932 11376 15960
rect 11422 15920 11428 15972
rect 11480 15960 11486 15972
rect 15470 15960 15476 15972
rect 11480 15932 15476 15960
rect 11480 15920 11486 15932
rect 15470 15920 15476 15932
rect 15528 15920 15534 15972
rect 9858 15852 9864 15904
rect 9916 15852 9922 15904
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11790 15892 11796 15904
rect 11112 15864 11796 15892
rect 11112 15852 11118 15864
rect 11790 15852 11796 15864
rect 11848 15892 11854 15904
rect 12253 15895 12311 15901
rect 12253 15892 12265 15895
rect 11848 15864 12265 15892
rect 11848 15852 11854 15864
rect 12253 15861 12265 15864
rect 12299 15861 12311 15895
rect 12253 15855 12311 15861
rect 13449 15895 13507 15901
rect 13449 15861 13461 15895
rect 13495 15892 13507 15895
rect 14642 15892 14648 15904
rect 13495 15864 14648 15892
rect 13495 15861 13507 15864
rect 13449 15855 13507 15861
rect 14642 15852 14648 15864
rect 14700 15852 14706 15904
rect 15838 15852 15844 15904
rect 15896 15892 15902 15904
rect 17954 15892 17960 15904
rect 15896 15864 17960 15892
rect 15896 15852 15902 15864
rect 17954 15852 17960 15864
rect 18012 15852 18018 15904
rect 1104 15802 18860 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 6950 15802
rect 7002 15750 7014 15802
rect 7066 15750 7078 15802
rect 7130 15750 7142 15802
rect 7194 15750 7206 15802
rect 7258 15750 11950 15802
rect 12002 15750 12014 15802
rect 12066 15750 12078 15802
rect 12130 15750 12142 15802
rect 12194 15750 12206 15802
rect 12258 15750 16950 15802
rect 17002 15750 17014 15802
rect 17066 15750 17078 15802
rect 17130 15750 17142 15802
rect 17194 15750 17206 15802
rect 17258 15750 18860 15802
rect 1104 15728 18860 15750
rect 10962 15648 10968 15700
rect 11020 15688 11026 15700
rect 11422 15688 11428 15700
rect 11020 15660 11428 15688
rect 11020 15648 11026 15660
rect 11422 15648 11428 15660
rect 11480 15648 11486 15700
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 14185 15691 14243 15697
rect 14185 15688 14197 15691
rect 14148 15660 14197 15688
rect 14148 15648 14154 15660
rect 14185 15657 14197 15660
rect 14231 15688 14243 15691
rect 14921 15691 14979 15697
rect 14921 15688 14933 15691
rect 14231 15660 14933 15688
rect 14231 15657 14243 15660
rect 14185 15651 14243 15657
rect 14921 15657 14933 15660
rect 14967 15657 14979 15691
rect 14921 15651 14979 15657
rect 5718 15580 5724 15632
rect 5776 15620 5782 15632
rect 5776 15592 17356 15620
rect 5776 15580 5782 15592
rect 2406 15512 2412 15564
rect 2464 15552 2470 15564
rect 2464 15524 8156 15552
rect 2464 15512 2470 15524
rect 6638 15444 6644 15496
rect 6696 15444 6702 15496
rect 8128 15493 8156 15524
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 10505 15555 10563 15561
rect 10505 15552 10517 15555
rect 8536 15524 10517 15552
rect 8536 15512 8542 15524
rect 10505 15521 10517 15524
rect 10551 15552 10563 15555
rect 10686 15552 10692 15564
rect 10551 15524 10692 15552
rect 10551 15521 10563 15524
rect 10505 15515 10563 15521
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 10962 15512 10968 15564
rect 11020 15512 11026 15564
rect 13538 15512 13544 15564
rect 13596 15512 13602 15564
rect 13722 15512 13728 15564
rect 13780 15552 13786 15564
rect 17328 15561 17356 15592
rect 17313 15555 17371 15561
rect 13780 15524 17264 15552
rect 13780 15512 13786 15524
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15453 6791 15487
rect 6733 15447 6791 15453
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 2958 15376 2964 15428
rect 3016 15416 3022 15428
rect 6748 15416 6776 15447
rect 8294 15444 8300 15496
rect 8352 15444 8358 15496
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 10468 15456 10609 15484
rect 10468 15444 10474 15456
rect 10597 15453 10609 15456
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 13170 15444 13176 15496
rect 13228 15444 13234 15496
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 14918 15484 14924 15496
rect 14507 15456 14924 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 14918 15444 14924 15456
rect 14976 15444 14982 15496
rect 15470 15444 15476 15496
rect 15528 15444 15534 15496
rect 16574 15444 16580 15496
rect 16632 15484 16638 15496
rect 16761 15487 16819 15493
rect 16761 15484 16773 15487
rect 16632 15456 16773 15484
rect 16632 15444 16638 15456
rect 16761 15453 16773 15456
rect 16807 15453 16819 15487
rect 16761 15447 16819 15453
rect 17126 15444 17132 15496
rect 17184 15444 17190 15496
rect 17236 15484 17264 15524
rect 17313 15521 17325 15555
rect 17359 15521 17371 15555
rect 18417 15555 18475 15561
rect 18417 15552 18429 15555
rect 17313 15515 17371 15521
rect 17420 15524 18429 15552
rect 17420 15484 17448 15524
rect 18417 15521 18429 15524
rect 18463 15521 18475 15555
rect 18417 15515 18475 15521
rect 17236 15456 17448 15484
rect 17957 15487 18015 15493
rect 17957 15453 17969 15487
rect 18003 15484 18015 15487
rect 18046 15484 18052 15496
rect 18003 15456 18052 15484
rect 18003 15453 18015 15456
rect 17957 15447 18015 15453
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 18233 15487 18291 15493
rect 18233 15484 18245 15487
rect 18196 15456 18245 15484
rect 18196 15444 18202 15456
rect 18233 15453 18245 15456
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 12894 15416 12900 15428
rect 3016 15388 6776 15416
rect 6840 15388 12900 15416
rect 3016 15376 3022 15388
rect 5810 15308 5816 15360
rect 5868 15348 5874 15360
rect 6089 15351 6147 15357
rect 6089 15348 6101 15351
rect 5868 15320 6101 15348
rect 5868 15308 5874 15320
rect 6089 15317 6101 15320
rect 6135 15317 6147 15351
rect 6089 15311 6147 15317
rect 6362 15308 6368 15360
rect 6420 15348 6426 15360
rect 6840 15348 6868 15388
rect 12894 15376 12900 15388
rect 12952 15376 12958 15428
rect 12989 15419 13047 15425
rect 12989 15385 13001 15419
rect 13035 15416 13047 15419
rect 13262 15416 13268 15428
rect 13035 15388 13268 15416
rect 13035 15385 13047 15388
rect 12989 15379 13047 15385
rect 13262 15376 13268 15388
rect 13320 15376 13326 15428
rect 15105 15419 15163 15425
rect 15105 15416 15117 15419
rect 13740 15388 15117 15416
rect 6420 15320 6868 15348
rect 6420 15308 6426 15320
rect 8110 15308 8116 15360
rect 8168 15348 8174 15360
rect 8205 15351 8263 15357
rect 8205 15348 8217 15351
rect 8168 15320 8217 15348
rect 8168 15308 8174 15320
rect 8205 15317 8217 15320
rect 8251 15317 8263 15351
rect 8205 15311 8263 15317
rect 9030 15308 9036 15360
rect 9088 15348 9094 15360
rect 13740 15348 13768 15388
rect 15105 15385 15117 15388
rect 15151 15385 15163 15419
rect 15105 15379 15163 15385
rect 15289 15419 15347 15425
rect 15289 15385 15301 15419
rect 15335 15416 15347 15419
rect 15378 15416 15384 15428
rect 15335 15388 15384 15416
rect 15335 15385 15347 15388
rect 15289 15379 15347 15385
rect 15378 15376 15384 15388
rect 15436 15376 15442 15428
rect 16850 15376 16856 15428
rect 16908 15376 16914 15428
rect 18690 15416 18696 15428
rect 18064 15388 18696 15416
rect 9088 15320 13768 15348
rect 14645 15351 14703 15357
rect 9088 15308 9094 15320
rect 14645 15317 14657 15351
rect 14691 15348 14703 15351
rect 17954 15348 17960 15360
rect 14691 15320 17960 15348
rect 14691 15317 14703 15320
rect 14645 15311 14703 15317
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 18064 15357 18092 15388
rect 18690 15376 18696 15388
rect 18748 15376 18754 15428
rect 18049 15351 18107 15357
rect 18049 15317 18061 15351
rect 18095 15317 18107 15351
rect 18049 15311 18107 15317
rect 1104 15258 18860 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 7610 15258
rect 7662 15206 7674 15258
rect 7726 15206 7738 15258
rect 7790 15206 7802 15258
rect 7854 15206 7866 15258
rect 7918 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 17610 15258
rect 17662 15206 17674 15258
rect 17726 15206 17738 15258
rect 17790 15206 17802 15258
rect 17854 15206 17866 15258
rect 17918 15206 18860 15258
rect 1104 15184 18860 15206
rect 3878 15104 3884 15156
rect 3936 15144 3942 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 3936 15116 8217 15144
rect 3936 15104 3942 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8205 15107 8263 15113
rect 8938 15104 8944 15156
rect 8996 15144 9002 15156
rect 9674 15144 9680 15156
rect 8996 15116 9680 15144
rect 8996 15104 9002 15116
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 9968 15116 10456 15144
rect 5534 15076 5540 15088
rect 2746 15048 5540 15076
rect 842 14968 848 15020
rect 900 15008 906 15020
rect 1489 15011 1547 15017
rect 1489 15008 1501 15011
rect 900 14980 1501 15008
rect 900 14968 906 14980
rect 1489 14977 1501 14980
rect 1535 14977 1547 15011
rect 1489 14971 1547 14977
rect 1673 14875 1731 14881
rect 1673 14841 1685 14875
rect 1719 14872 1731 14875
rect 2746 14872 2774 15048
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 5644 15048 8156 15076
rect 3329 15011 3387 15017
rect 3329 14977 3341 15011
rect 3375 14977 3387 15011
rect 3329 14971 3387 14977
rect 3344 14940 3372 14971
rect 3510 14968 3516 15020
rect 3568 14968 3574 15020
rect 5644 15017 5672 15048
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 14977 5687 15011
rect 5629 14971 5687 14977
rect 5721 15011 5779 15017
rect 5721 14977 5733 15011
rect 5767 15008 5779 15011
rect 6638 15008 6644 15020
rect 5767 14980 6644 15008
rect 5767 14977 5779 14980
rect 5721 14971 5779 14977
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 7650 14968 7656 15020
rect 7708 14968 7714 15020
rect 8128 15017 8156 15048
rect 8570 15036 8576 15088
rect 8628 15076 8634 15088
rect 9398 15076 9404 15088
rect 8628 15048 9404 15076
rect 8628 15036 8634 15048
rect 9398 15036 9404 15048
rect 9456 15076 9462 15088
rect 9968 15076 9996 15116
rect 10428 15076 10456 15116
rect 10686 15104 10692 15156
rect 10744 15144 10750 15156
rect 10744 15116 13952 15144
rect 10744 15104 10750 15116
rect 9456 15048 9996 15076
rect 10060 15048 10364 15076
rect 10428 15048 11560 15076
rect 9456 15036 9462 15048
rect 7929 15011 7987 15017
rect 7929 14977 7941 15011
rect 7975 14977 7987 15011
rect 7929 14971 7987 14977
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 15008 8171 15011
rect 8202 15008 8208 15020
rect 8159 14980 8208 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 3344 14912 5948 14940
rect 1719 14844 2774 14872
rect 1719 14841 1731 14844
rect 1673 14835 1731 14841
rect 3237 14807 3295 14813
rect 3237 14773 3249 14807
rect 3283 14804 3295 14807
rect 3418 14804 3424 14816
rect 3283 14776 3424 14804
rect 3283 14773 3295 14776
rect 3237 14767 3295 14773
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 5920 14813 5948 14912
rect 7466 14900 7472 14952
rect 7524 14940 7530 14952
rect 7944 14940 7972 14971
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 15008 8355 15011
rect 8343 14980 9356 15008
rect 8343 14977 8355 14980
rect 8297 14971 8355 14977
rect 7524 14912 7972 14940
rect 7524 14900 7530 14912
rect 6730 14832 6736 14884
rect 6788 14872 6794 14884
rect 7745 14875 7803 14881
rect 7745 14872 7757 14875
rect 6788 14844 7757 14872
rect 6788 14832 6794 14844
rect 7745 14841 7757 14844
rect 7791 14841 7803 14875
rect 7745 14835 7803 14841
rect 7837 14875 7895 14881
rect 7837 14841 7849 14875
rect 7883 14872 7895 14875
rect 8018 14872 8024 14884
rect 7883 14844 8024 14872
rect 7883 14841 7895 14844
rect 7837 14835 7895 14841
rect 5905 14807 5963 14813
rect 5905 14773 5917 14807
rect 5951 14804 5963 14807
rect 6086 14804 6092 14816
rect 5951 14776 6092 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 6086 14764 6092 14776
rect 6144 14764 6150 14816
rect 7469 14807 7527 14813
rect 7469 14773 7481 14807
rect 7515 14804 7527 14807
rect 7558 14804 7564 14816
rect 7515 14776 7564 14804
rect 7515 14773 7527 14776
rect 7469 14767 7527 14773
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 7760 14804 7788 14835
rect 8018 14832 8024 14844
rect 8076 14832 8082 14884
rect 8662 14832 8668 14884
rect 8720 14872 8726 14884
rect 9125 14875 9183 14881
rect 9125 14872 9137 14875
rect 8720 14844 9137 14872
rect 8720 14832 8726 14844
rect 9125 14841 9137 14844
rect 9171 14841 9183 14875
rect 9328 14872 9356 14980
rect 9674 14968 9680 15020
rect 9732 14968 9738 15020
rect 9953 15014 10011 15017
rect 10060 15014 10088 15048
rect 9953 15011 10088 15014
rect 9953 14977 9965 15011
rect 9999 14986 10088 15011
rect 10336 15008 10364 15048
rect 10594 15008 10600 15020
rect 9999 14977 10011 14986
rect 10336 14980 10600 15008
rect 9953 14971 10011 14977
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 11532 15008 11560 15048
rect 12618 15036 12624 15088
rect 12676 15076 12682 15088
rect 13722 15076 13728 15088
rect 12676 15048 13728 15076
rect 12676 15036 12682 15048
rect 13722 15036 13728 15048
rect 13780 15036 13786 15088
rect 11606 15008 11612 15020
rect 11532 14980 11612 15008
rect 11606 14968 11612 14980
rect 11664 15008 11670 15020
rect 13924 15017 13952 15116
rect 17862 15104 17868 15156
rect 17920 15144 17926 15156
rect 18322 15144 18328 15156
rect 17920 15116 18328 15144
rect 17920 15104 17926 15116
rect 18322 15104 18328 15116
rect 18380 15104 18386 15156
rect 17126 15036 17132 15088
rect 17184 15076 17190 15088
rect 17954 15076 17960 15088
rect 17184 15048 17960 15076
rect 17184 15036 17190 15048
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 11664 14980 13369 15008
rect 11664 14968 11670 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 13909 15011 13967 15017
rect 13909 14977 13921 15011
rect 13955 14977 13967 15011
rect 13909 14971 13967 14977
rect 14182 14968 14188 15020
rect 14240 15008 14246 15020
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 14240 14980 14473 15008
rect 14240 14968 14246 14980
rect 14461 14977 14473 14980
rect 14507 15008 14519 15011
rect 14550 15008 14556 15020
rect 14507 14980 14556 15008
rect 14507 14977 14519 14980
rect 14461 14971 14519 14977
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 16114 14968 16120 15020
rect 16172 15008 16178 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16172 14980 16865 15008
rect 16172 14968 16178 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 16945 15011 17003 15017
rect 16945 14977 16957 15011
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17267 14980 17540 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 9398 14900 9404 14952
rect 9456 14900 9462 14952
rect 9766 14900 9772 14952
rect 9824 14940 9830 14952
rect 9861 14943 9919 14949
rect 9861 14940 9873 14943
rect 9824 14912 9873 14940
rect 9824 14900 9830 14912
rect 9861 14909 9873 14912
rect 9907 14909 9919 14943
rect 9861 14903 9919 14909
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14909 10103 14943
rect 10045 14903 10103 14909
rect 9674 14872 9680 14884
rect 9328 14844 9680 14872
rect 9125 14835 9183 14841
rect 9674 14832 9680 14844
rect 9732 14832 9738 14884
rect 10060 14872 10088 14903
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10192 14912 10236 14940
rect 10192 14900 10198 14912
rect 12894 14900 12900 14952
rect 12952 14940 12958 14952
rect 14090 14940 14096 14952
rect 12952 14912 14096 14940
rect 12952 14900 12958 14912
rect 14090 14900 14096 14912
rect 14148 14900 14154 14952
rect 14366 14900 14372 14952
rect 14424 14940 14430 14952
rect 15197 14943 15255 14949
rect 15197 14940 15209 14943
rect 14424 14912 15209 14940
rect 14424 14900 14430 14912
rect 15197 14909 15209 14912
rect 15243 14909 15255 14943
rect 15197 14903 15255 14909
rect 16758 14900 16764 14952
rect 16816 14940 16822 14952
rect 16960 14940 16988 14971
rect 17512 14952 17540 14980
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 18598 15008 18604 15020
rect 18380 14980 18604 15008
rect 18380 14968 18386 14980
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 16816 14912 16988 14940
rect 16816 14900 16822 14912
rect 17494 14900 17500 14952
rect 17552 14900 17558 14952
rect 10502 14872 10508 14884
rect 10060 14844 10508 14872
rect 10502 14832 10508 14844
rect 10560 14832 10566 14884
rect 14826 14832 14832 14884
rect 14884 14832 14890 14884
rect 8938 14804 8944 14816
rect 7760 14776 8944 14804
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 9490 14764 9496 14816
rect 9548 14764 9554 14816
rect 10321 14807 10379 14813
rect 10321 14773 10333 14807
rect 10367 14804 10379 14807
rect 13538 14804 13544 14816
rect 10367 14776 13544 14804
rect 10367 14773 10379 14776
rect 10321 14767 10379 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 13725 14807 13783 14813
rect 13725 14773 13737 14807
rect 13771 14804 13783 14807
rect 14458 14804 14464 14816
rect 13771 14776 14464 14804
rect 13771 14773 13783 14776
rect 13725 14767 13783 14773
rect 14458 14764 14464 14776
rect 14516 14764 14522 14816
rect 14734 14764 14740 14816
rect 14792 14764 14798 14816
rect 16574 14764 16580 14816
rect 16632 14804 16638 14816
rect 16669 14807 16727 14813
rect 16669 14804 16681 14807
rect 16632 14776 16681 14804
rect 16632 14764 16638 14776
rect 16669 14773 16681 14776
rect 16715 14773 16727 14807
rect 16669 14767 16727 14773
rect 17129 14807 17187 14813
rect 17129 14773 17141 14807
rect 17175 14804 17187 14807
rect 18874 14804 18880 14816
rect 17175 14776 18880 14804
rect 17175 14773 17187 14776
rect 17129 14767 17187 14773
rect 18874 14764 18880 14776
rect 18932 14764 18938 14816
rect 1104 14714 18860 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 6950 14714
rect 7002 14662 7014 14714
rect 7066 14662 7078 14714
rect 7130 14662 7142 14714
rect 7194 14662 7206 14714
rect 7258 14662 11950 14714
rect 12002 14662 12014 14714
rect 12066 14662 12078 14714
rect 12130 14662 12142 14714
rect 12194 14662 12206 14714
rect 12258 14662 16950 14714
rect 17002 14662 17014 14714
rect 17066 14662 17078 14714
rect 17130 14662 17142 14714
rect 17194 14662 17206 14714
rect 17258 14662 18860 14714
rect 1104 14640 18860 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 7650 14600 7656 14612
rect 1912 14572 7656 14600
rect 1912 14560 1918 14572
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 9674 14600 9680 14612
rect 8312 14572 9680 14600
rect 8312 14544 8340 14572
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 10134 14560 10140 14612
rect 10192 14600 10198 14612
rect 12618 14600 12624 14612
rect 10192 14572 12624 14600
rect 10192 14560 10198 14572
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 14918 14600 14924 14612
rect 13596 14572 14924 14600
rect 13596 14560 13602 14572
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 8294 14532 8300 14544
rect 4212 14504 8300 14532
rect 4212 14492 4218 14504
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 8570 14492 8576 14544
rect 8628 14532 8634 14544
rect 9401 14535 9459 14541
rect 9401 14532 9413 14535
rect 8628 14504 9413 14532
rect 8628 14492 8634 14504
rect 9401 14501 9413 14504
rect 9447 14532 9459 14535
rect 12894 14532 12900 14544
rect 9447 14504 12900 14532
rect 9447 14501 9459 14504
rect 9401 14495 9459 14501
rect 12894 14492 12900 14504
rect 12952 14492 12958 14544
rect 13078 14492 13084 14544
rect 13136 14532 13142 14544
rect 13446 14532 13452 14544
rect 13136 14504 13452 14532
rect 13136 14492 13142 14504
rect 13446 14492 13452 14504
rect 13504 14492 13510 14544
rect 14090 14492 14096 14544
rect 14148 14532 14154 14544
rect 16669 14535 16727 14541
rect 16669 14532 16681 14535
rect 14148 14504 16681 14532
rect 14148 14492 14154 14504
rect 16669 14501 16681 14504
rect 16715 14501 16727 14535
rect 16669 14495 16727 14501
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 7616 14453 10180 14464
rect 10226 14453 10232 14476
rect 7616 14436 10232 14453
rect 7616 14424 7622 14436
rect 10152 14425 10232 14436
rect 10226 14424 10232 14425
rect 10284 14424 10290 14476
rect 10321 14467 10379 14473
rect 10321 14433 10333 14467
rect 10367 14464 10379 14467
rect 10502 14464 10508 14476
rect 10367 14436 10508 14464
rect 10367 14433 10379 14436
rect 10321 14427 10379 14433
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 13354 14424 13360 14476
rect 13412 14464 13418 14476
rect 15746 14464 15752 14476
rect 13412 14436 15752 14464
rect 13412 14424 13418 14436
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 18414 14464 18420 14476
rect 16868 14436 18420 14464
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 16868 14405 16896 14436
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 10045 14399 10103 14405
rect 10045 14396 10057 14399
rect 8168 14368 10057 14396
rect 8168 14356 8174 14368
rect 10045 14365 10057 14368
rect 10091 14365 10103 14399
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 10045 14359 10103 14365
rect 10244 14368 14657 14396
rect 5902 14288 5908 14340
rect 5960 14328 5966 14340
rect 9125 14331 9183 14337
rect 9125 14328 9137 14331
rect 5960 14300 9137 14328
rect 5960 14288 5966 14300
rect 9125 14297 9137 14300
rect 9171 14297 9183 14331
rect 10244 14328 10272 14368
rect 14645 14365 14657 14368
rect 14691 14365 14703 14399
rect 14829 14399 14887 14405
rect 14829 14396 14841 14399
rect 14645 14359 14703 14365
rect 14752 14368 14841 14396
rect 9125 14291 9183 14297
rect 9232 14300 10272 14328
rect 10321 14331 10379 14337
rect 8018 14220 8024 14272
rect 8076 14260 8082 14272
rect 9232 14260 9260 14300
rect 10321 14297 10333 14331
rect 10367 14328 10379 14331
rect 11698 14328 11704 14340
rect 10367 14300 11704 14328
rect 10367 14297 10379 14300
rect 10321 14291 10379 14297
rect 11698 14288 11704 14300
rect 11756 14288 11762 14340
rect 8076 14232 9260 14260
rect 8076 14220 8082 14232
rect 9582 14220 9588 14272
rect 9640 14220 9646 14272
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 14752 14260 14780 14368
rect 14829 14365 14841 14368
rect 14875 14365 14887 14399
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 14829 14359 14887 14365
rect 15212 14368 16865 14396
rect 11020 14232 14780 14260
rect 11020 14220 11026 14232
rect 14918 14220 14924 14272
rect 14976 14260 14982 14272
rect 15212 14260 15240 14368
rect 16853 14365 16865 14368
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 17129 14399 17187 14405
rect 17129 14365 17141 14399
rect 17175 14396 17187 14399
rect 17862 14396 17868 14408
rect 17175 14368 17868 14396
rect 17175 14365 17187 14368
rect 17129 14359 17187 14365
rect 16758 14288 16764 14340
rect 16816 14328 16822 14340
rect 17144 14328 17172 14359
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 16816 14300 17172 14328
rect 16816 14288 16822 14300
rect 14976 14232 15240 14260
rect 14976 14220 14982 14232
rect 15654 14220 15660 14272
rect 15712 14220 15718 14272
rect 17034 14220 17040 14272
rect 17092 14260 17098 14272
rect 17402 14260 17408 14272
rect 17092 14232 17408 14260
rect 17092 14220 17098 14232
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 1104 14170 18860 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 7610 14170
rect 7662 14118 7674 14170
rect 7726 14118 7738 14170
rect 7790 14118 7802 14170
rect 7854 14118 7866 14170
rect 7918 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 17610 14170
rect 17662 14118 17674 14170
rect 17726 14118 17738 14170
rect 17790 14118 17802 14170
rect 17854 14118 17866 14170
rect 17918 14118 18860 14170
rect 1104 14096 18860 14118
rect 7558 14016 7564 14068
rect 7616 14056 7622 14068
rect 8202 14056 8208 14068
rect 7616 14028 8208 14056
rect 7616 14016 7622 14028
rect 8202 14016 8208 14028
rect 8260 14016 8266 14068
rect 9217 14059 9275 14065
rect 8772 14028 9168 14056
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 8662 13988 8668 14000
rect 8076 13960 8668 13988
rect 8076 13948 8082 13960
rect 8662 13948 8668 13960
rect 8720 13948 8726 14000
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 5258 13880 5264 13932
rect 5316 13920 5322 13932
rect 8772 13929 8800 14028
rect 9140 13988 9168 14028
rect 9217 14025 9229 14059
rect 9263 14056 9275 14059
rect 9306 14056 9312 14068
rect 9263 14028 9312 14056
rect 9263 14025 9275 14028
rect 9217 14019 9275 14025
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 9398 14016 9404 14068
rect 9456 14056 9462 14068
rect 9582 14056 9588 14068
rect 9456 14028 9588 14056
rect 9456 14016 9462 14028
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 10226 14016 10232 14068
rect 10284 14056 10290 14068
rect 10284 14028 14688 14056
rect 10284 14016 10290 14028
rect 12342 13988 12348 14000
rect 9140 13960 12348 13988
rect 12342 13948 12348 13960
rect 12400 13948 12406 14000
rect 12437 13991 12495 13997
rect 12437 13957 12449 13991
rect 12483 13988 12495 13991
rect 12526 13988 12532 14000
rect 12483 13960 12532 13988
rect 12483 13957 12495 13960
rect 12437 13951 12495 13957
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 12621 13991 12679 13997
rect 12621 13957 12633 13991
rect 12667 13988 12679 13991
rect 13354 13988 13360 14000
rect 12667 13960 13360 13988
rect 12667 13957 12679 13960
rect 12621 13951 12679 13957
rect 13354 13948 13360 13960
rect 13412 13948 13418 14000
rect 8757 13923 8815 13929
rect 5316 13892 7880 13920
rect 5316 13880 5322 13892
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 6178 13852 6184 13864
rect 3476 13824 6184 13852
rect 3476 13812 3482 13824
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 7852 13852 7880 13892
rect 8757 13889 8769 13923
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 9030 13880 9036 13932
rect 9088 13880 9094 13932
rect 9122 13880 9128 13932
rect 9180 13920 9186 13932
rect 10042 13920 10048 13932
rect 9180 13892 10048 13920
rect 9180 13880 9186 13892
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13920 13967 13923
rect 14366 13920 14372 13932
rect 13955 13892 14372 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 14550 13880 14556 13932
rect 14608 13880 14614 13932
rect 14660 13929 14688 14028
rect 18414 14016 18420 14068
rect 18472 14016 18478 14068
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 14826 13880 14832 13932
rect 14884 13880 14890 13932
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 18233 13923 18291 13929
rect 18233 13920 18245 13923
rect 15344 13892 18245 13920
rect 15344 13880 15350 13892
rect 18233 13889 18245 13892
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 8662 13852 8668 13864
rect 7852 13824 8668 13852
rect 8662 13812 8668 13824
rect 8720 13852 8726 13864
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8720 13824 8861 13852
rect 8720 13812 8726 13824
rect 8849 13821 8861 13824
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 8941 13855 8999 13861
rect 8941 13821 8953 13855
rect 8987 13852 8999 13855
rect 11422 13852 11428 13864
rect 8987 13824 11428 13852
rect 8987 13821 8999 13824
rect 8941 13815 8999 13821
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 13630 13812 13636 13864
rect 13688 13812 13694 13864
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 14918 13852 14924 13864
rect 14056 13824 14924 13852
rect 14056 13812 14062 13824
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 1670 13744 1676 13796
rect 1728 13784 1734 13796
rect 6914 13784 6920 13796
rect 1728 13756 6920 13784
rect 1728 13744 1734 13756
rect 6914 13744 6920 13756
rect 6972 13784 6978 13796
rect 8202 13784 8208 13796
rect 6972 13756 8208 13784
rect 6972 13744 6978 13756
rect 8202 13744 8208 13756
rect 8260 13744 8266 13796
rect 8386 13744 8392 13796
rect 8444 13784 8450 13796
rect 15013 13787 15071 13793
rect 15013 13784 15025 13787
rect 8444 13756 15025 13784
rect 8444 13744 8450 13756
rect 15013 13753 15025 13756
rect 15059 13753 15071 13787
rect 15013 13747 15071 13753
rect 15102 13744 15108 13796
rect 15160 13784 15166 13796
rect 15562 13784 15568 13796
rect 15160 13756 15568 13784
rect 15160 13744 15166 13756
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 1581 13719 1639 13725
rect 1581 13685 1593 13719
rect 1627 13716 1639 13719
rect 1762 13716 1768 13728
rect 1627 13688 1768 13716
rect 1627 13685 1639 13688
rect 1581 13679 1639 13685
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 6454 13676 6460 13728
rect 6512 13716 6518 13728
rect 8110 13716 8116 13728
rect 6512 13688 8116 13716
rect 6512 13676 6518 13688
rect 8110 13676 8116 13688
rect 8168 13676 8174 13728
rect 9030 13676 9036 13728
rect 9088 13716 9094 13728
rect 11514 13716 11520 13728
rect 9088 13688 11520 13716
rect 9088 13676 9094 13688
rect 11514 13676 11520 13688
rect 11572 13716 11578 13728
rect 12253 13719 12311 13725
rect 12253 13716 12265 13719
rect 11572 13688 12265 13716
rect 11572 13676 11578 13688
rect 12253 13685 12265 13688
rect 12299 13685 12311 13719
rect 12253 13679 12311 13685
rect 12526 13676 12532 13728
rect 12584 13716 12590 13728
rect 13538 13716 13544 13728
rect 12584 13688 13544 13716
rect 12584 13676 12590 13688
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 13909 13719 13967 13725
rect 13909 13685 13921 13719
rect 13955 13716 13967 13719
rect 15470 13716 15476 13728
rect 13955 13688 15476 13716
rect 13955 13685 13967 13688
rect 13909 13679 13967 13685
rect 15470 13676 15476 13688
rect 15528 13716 15534 13728
rect 18138 13716 18144 13728
rect 15528 13688 18144 13716
rect 15528 13676 15534 13688
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 1104 13626 18860 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 11950 13626
rect 12002 13574 12014 13626
rect 12066 13574 12078 13626
rect 12130 13574 12142 13626
rect 12194 13574 12206 13626
rect 12258 13574 16950 13626
rect 17002 13574 17014 13626
rect 17066 13574 17078 13626
rect 17130 13574 17142 13626
rect 17194 13574 17206 13626
rect 17258 13574 18860 13626
rect 1104 13552 18860 13574
rect 6638 13472 6644 13524
rect 6696 13512 6702 13524
rect 7190 13512 7196 13524
rect 6696 13484 7196 13512
rect 6696 13472 6702 13484
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7926 13472 7932 13524
rect 7984 13512 7990 13524
rect 8110 13512 8116 13524
rect 7984 13484 8116 13512
rect 7984 13472 7990 13484
rect 8110 13472 8116 13484
rect 8168 13512 8174 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8168 13484 9045 13512
rect 8168 13472 8174 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 9033 13475 9091 13481
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 10100 13484 10916 13512
rect 10100 13472 10106 13484
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 8938 13444 8944 13456
rect 5592 13416 8944 13444
rect 5592 13404 5598 13416
rect 8938 13404 8944 13416
rect 8996 13444 9002 13456
rect 9313 13447 9371 13453
rect 9313 13444 9325 13447
rect 8996 13416 9325 13444
rect 8996 13404 9002 13416
rect 9313 13413 9325 13416
rect 9359 13413 9371 13447
rect 9313 13407 9371 13413
rect 9401 13447 9459 13453
rect 9401 13413 9413 13447
rect 9447 13444 9459 13447
rect 10778 13444 10784 13456
rect 9447 13416 10784 13444
rect 9447 13413 9459 13416
rect 9401 13407 9459 13413
rect 10778 13404 10784 13416
rect 10836 13404 10842 13456
rect 10888 13444 10916 13484
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 13538 13512 13544 13524
rect 13228 13484 13544 13512
rect 13228 13472 13234 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 17494 13512 17500 13524
rect 14200 13484 17500 13512
rect 13814 13444 13820 13456
rect 10888 13416 13820 13444
rect 13814 13404 13820 13416
rect 13872 13404 13878 13456
rect 3786 13336 3792 13388
rect 3844 13376 3850 13388
rect 6917 13379 6975 13385
rect 6917 13376 6929 13379
rect 3844 13348 6929 13376
rect 3844 13336 3850 13348
rect 6917 13345 6929 13348
rect 6963 13376 6975 13379
rect 10962 13376 10968 13388
rect 6963 13348 10968 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 11422 13336 11428 13388
rect 11480 13376 11486 13388
rect 12250 13376 12256 13388
rect 11480 13348 12256 13376
rect 11480 13336 11486 13348
rect 12250 13336 12256 13348
rect 12308 13376 12314 13388
rect 12805 13379 12863 13385
rect 12805 13376 12817 13379
rect 12308 13348 12817 13376
rect 12308 13336 12314 13348
rect 12805 13345 12817 13348
rect 12851 13345 12863 13379
rect 12805 13339 12863 13345
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13376 13047 13379
rect 13354 13376 13360 13388
rect 13035 13348 13360 13376
rect 13035 13345 13047 13348
rect 12989 13339 13047 13345
rect 13354 13336 13360 13348
rect 13412 13376 13418 13388
rect 14090 13376 14096 13388
rect 13412 13348 14096 13376
rect 13412 13336 13418 13348
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 2958 13268 2964 13320
rect 3016 13308 3022 13320
rect 3145 13311 3203 13317
rect 3145 13308 3157 13311
rect 3016 13280 3157 13308
rect 3016 13268 3022 13280
rect 3145 13277 3157 13280
rect 3191 13277 3203 13311
rect 3145 13271 3203 13277
rect 3326 13268 3332 13320
rect 3384 13268 3390 13320
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13308 3571 13311
rect 5718 13308 5724 13320
rect 3559 13280 5724 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 9030 13308 9036 13320
rect 7055 13280 9036 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 9214 13268 9220 13320
rect 9272 13268 9278 13320
rect 9398 13268 9404 13320
rect 9456 13308 9462 13320
rect 9493 13311 9551 13317
rect 9493 13308 9505 13311
rect 9456 13280 9505 13308
rect 9456 13268 9462 13280
rect 9493 13277 9505 13280
rect 9539 13277 9551 13311
rect 9493 13271 9551 13277
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 12526 13308 12532 13320
rect 9824 13280 12532 13308
rect 9824 13268 9830 13280
rect 12526 13268 12532 13280
rect 12584 13268 12590 13320
rect 12710 13268 12716 13320
rect 12768 13268 12774 13320
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13308 12955 13311
rect 13722 13308 13728 13320
rect 12943 13280 13728 13308
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 13722 13268 13728 13280
rect 13780 13308 13786 13320
rect 14200 13308 14228 13484
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 15194 13404 15200 13456
rect 15252 13444 15258 13456
rect 15252 13416 15976 13444
rect 15252 13404 15258 13416
rect 14737 13379 14795 13385
rect 14737 13345 14749 13379
rect 14783 13376 14795 13379
rect 15654 13376 15660 13388
rect 14783 13348 15660 13376
rect 14783 13345 14795 13348
rect 14737 13339 14795 13345
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 15948 13385 15976 13416
rect 15933 13379 15991 13385
rect 15933 13345 15945 13379
rect 15979 13376 15991 13379
rect 16206 13376 16212 13388
rect 15979 13348 16212 13376
rect 15979 13345 15991 13348
rect 15933 13339 15991 13345
rect 16206 13336 16212 13348
rect 16264 13336 16270 13388
rect 13780 13280 14228 13308
rect 13780 13268 13786 13280
rect 14550 13268 14556 13320
rect 14608 13268 14614 13320
rect 14826 13268 14832 13320
rect 14884 13308 14890 13320
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 14884 13280 15485 13308
rect 14884 13268 14890 13280
rect 15473 13277 15485 13280
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 15562 13268 15568 13320
rect 15620 13308 15626 13320
rect 16022 13308 16028 13320
rect 15620 13280 16028 13308
rect 15620 13268 15626 13280
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 3602 13200 3608 13252
rect 3660 13240 3666 13252
rect 3970 13240 3976 13252
rect 3660 13212 3976 13240
rect 3660 13200 3666 13212
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 9582 13200 9588 13252
rect 9640 13240 9646 13252
rect 14458 13240 14464 13252
rect 9640 13212 14464 13240
rect 9640 13200 9646 13212
rect 14458 13200 14464 13212
rect 14516 13240 14522 13252
rect 15105 13243 15163 13249
rect 15105 13240 15117 13243
rect 14516 13212 15117 13240
rect 14516 13200 14522 13212
rect 15105 13209 15117 13212
rect 15151 13209 15163 13243
rect 15105 13203 15163 13209
rect 4522 13132 4528 13184
rect 4580 13172 4586 13184
rect 8386 13172 8392 13184
rect 4580 13144 8392 13172
rect 4580 13132 4586 13144
rect 8386 13132 8392 13144
rect 8444 13172 8450 13184
rect 8754 13172 8760 13184
rect 8444 13144 8760 13172
rect 8444 13132 8450 13144
rect 8754 13132 8760 13144
rect 8812 13132 8818 13184
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 14090 13172 14096 13184
rect 11020 13144 14096 13172
rect 11020 13132 11026 13144
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 1104 13082 18860 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 7610 13082
rect 7662 13030 7674 13082
rect 7726 13030 7738 13082
rect 7790 13030 7802 13082
rect 7854 13030 7866 13082
rect 7918 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 17610 13082
rect 17662 13030 17674 13082
rect 17726 13030 17738 13082
rect 17790 13030 17802 13082
rect 17854 13030 17866 13082
rect 17918 13030 18860 13082
rect 1104 13008 18860 13030
rect 1486 12928 1492 12980
rect 1544 12968 1550 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 1544 12940 1593 12968
rect 1544 12928 1550 12940
rect 1581 12937 1593 12940
rect 1627 12968 1639 12971
rect 1854 12968 1860 12980
rect 1627 12940 1860 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 3053 12971 3111 12977
rect 3053 12937 3065 12971
rect 3099 12968 3111 12971
rect 5902 12968 5908 12980
rect 3099 12940 5908 12968
rect 3099 12937 3111 12940
rect 3053 12931 3111 12937
rect 5902 12928 5908 12940
rect 5960 12928 5966 12980
rect 7377 12971 7435 12977
rect 7377 12937 7389 12971
rect 7423 12968 7435 12971
rect 10318 12968 10324 12980
rect 7423 12940 10324 12968
rect 7423 12937 7435 12940
rect 7377 12931 7435 12937
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10410 12928 10416 12980
rect 10468 12968 10474 12980
rect 10505 12971 10563 12977
rect 10505 12968 10517 12971
rect 10468 12940 10517 12968
rect 10468 12928 10474 12940
rect 10505 12937 10517 12940
rect 10551 12968 10563 12971
rect 13078 12968 13084 12980
rect 10551 12940 13084 12968
rect 10551 12937 10563 12940
rect 10505 12931 10563 12937
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 13630 12968 13636 12980
rect 13320 12940 13636 12968
rect 13320 12928 13326 12940
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 14274 12928 14280 12980
rect 14332 12968 14338 12980
rect 14550 12968 14556 12980
rect 14332 12940 14556 12968
rect 14332 12928 14338 12940
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 6089 12903 6147 12909
rect 6089 12869 6101 12903
rect 6135 12900 6147 12903
rect 14366 12900 14372 12912
rect 6135 12872 14372 12900
rect 6135 12869 6147 12872
rect 6089 12863 6147 12869
rect 14366 12860 14372 12872
rect 14424 12900 14430 12912
rect 17494 12900 17500 12912
rect 14424 12872 17500 12900
rect 14424 12860 14430 12872
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 842 12792 848 12844
rect 900 12832 906 12844
rect 1397 12835 1455 12841
rect 1397 12832 1409 12835
rect 900 12804 1409 12832
rect 900 12792 906 12804
rect 1397 12801 1409 12804
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12832 3387 12835
rect 3418 12832 3424 12844
rect 3375 12804 3424 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 3786 12792 3792 12844
rect 3844 12792 3850 12844
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12832 4215 12835
rect 4430 12832 4436 12844
rect 4203 12804 4436 12832
rect 4203 12801 4215 12804
rect 4157 12795 4215 12801
rect 4430 12792 4436 12804
rect 4488 12792 4494 12844
rect 4522 12792 4528 12844
rect 4580 12792 4586 12844
rect 4890 12792 4896 12844
rect 4948 12792 4954 12844
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 5626 12832 5632 12844
rect 5491 12804 5632 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 5718 12792 5724 12844
rect 5776 12792 5782 12844
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12832 7343 12835
rect 7466 12832 7472 12844
rect 7331 12804 7472 12832
rect 7331 12801 7343 12804
rect 7285 12795 7343 12801
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12832 7803 12835
rect 7834 12832 7840 12844
rect 7791 12804 7840 12832
rect 7791 12801 7803 12804
rect 7745 12795 7803 12801
rect 7834 12792 7840 12804
rect 7892 12792 7898 12844
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12832 8171 12835
rect 8202 12832 8208 12844
rect 8159 12804 8208 12832
rect 8159 12801 8171 12804
rect 8113 12795 8171 12801
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 8294 12792 8300 12844
rect 8352 12792 8358 12844
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 9582 12832 9588 12844
rect 8904 12804 9588 12832
rect 8904 12792 8910 12804
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 10318 12792 10324 12844
rect 10376 12832 10382 12844
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 10376 12804 10425 12832
rect 10376 12792 10382 12804
rect 10413 12801 10425 12804
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 7653 12767 7711 12773
rect 6871 12736 7604 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 5718 12656 5724 12708
rect 5776 12656 5782 12708
rect 7193 12699 7251 12705
rect 7193 12665 7205 12699
rect 7239 12696 7251 12699
rect 7282 12696 7288 12708
rect 7239 12668 7288 12696
rect 7239 12665 7251 12668
rect 7193 12659 7251 12665
rect 7282 12656 7288 12668
rect 7340 12656 7346 12708
rect 7576 12696 7604 12736
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 8754 12764 8760 12776
rect 7699 12736 8760 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 10428 12764 10456 12795
rect 10502 12792 10508 12844
rect 10560 12832 10566 12844
rect 10686 12832 10692 12844
rect 10560 12804 10692 12832
rect 10560 12792 10566 12804
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 11790 12792 11796 12844
rect 11848 12832 11854 12844
rect 12250 12832 12256 12844
rect 11848 12804 12256 12832
rect 11848 12792 11854 12804
rect 12250 12792 12256 12804
rect 12308 12832 12314 12844
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 12308 12804 13737 12832
rect 12308 12792 12314 12804
rect 13725 12801 13737 12804
rect 13771 12801 13783 12835
rect 13725 12795 13783 12801
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 14918 12832 14924 12844
rect 13872 12804 14924 12832
rect 13872 12792 13878 12804
rect 14918 12792 14924 12804
rect 14976 12792 14982 12844
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 10428 12736 13645 12764
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12764 13967 12767
rect 16758 12764 16764 12776
rect 13955 12736 16764 12764
rect 13955 12733 13967 12736
rect 13909 12727 13967 12733
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 7926 12696 7932 12708
rect 7576 12668 7932 12696
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 8386 12656 8392 12708
rect 8444 12696 8450 12708
rect 11422 12696 11428 12708
rect 8444 12668 11428 12696
rect 8444 12656 8450 12668
rect 11422 12656 11428 12668
rect 11480 12656 11486 12708
rect 12986 12696 12992 12708
rect 12406 12668 12992 12696
rect 5736 12628 5764 12656
rect 7374 12628 7380 12640
rect 5736 12600 7380 12628
rect 7374 12588 7380 12600
rect 7432 12588 7438 12640
rect 7742 12588 7748 12640
rect 7800 12588 7806 12640
rect 8202 12588 8208 12640
rect 8260 12588 8266 12640
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 12406 12628 12434 12668
rect 12986 12656 12992 12668
rect 13044 12696 13050 12708
rect 14274 12696 14280 12708
rect 13044 12668 14280 12696
rect 13044 12656 13050 12668
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 8720 12600 12434 12628
rect 8720 12588 8726 12600
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 13449 12631 13507 12637
rect 13449 12628 13461 12631
rect 12584 12600 13461 12628
rect 12584 12588 12590 12600
rect 13449 12597 13461 12600
rect 13495 12597 13507 12631
rect 13449 12591 13507 12597
rect 1104 12538 18860 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 11950 12538
rect 12002 12486 12014 12538
rect 12066 12486 12078 12538
rect 12130 12486 12142 12538
rect 12194 12486 12206 12538
rect 12258 12486 16950 12538
rect 17002 12486 17014 12538
rect 17066 12486 17078 12538
rect 17130 12486 17142 12538
rect 17194 12486 17206 12538
rect 17258 12486 18860 12538
rect 1104 12464 18860 12486
rect 1578 12384 1584 12436
rect 1636 12424 1642 12436
rect 1636 12396 7420 12424
rect 1636 12384 1642 12396
rect 1762 12316 1768 12368
rect 1820 12356 1826 12368
rect 6730 12356 6736 12368
rect 1820 12328 6736 12356
rect 1820 12316 1826 12328
rect 6730 12316 6736 12328
rect 6788 12356 6794 12368
rect 7392 12356 7420 12396
rect 8110 12384 8116 12436
rect 8168 12424 8174 12436
rect 9585 12427 9643 12433
rect 8168 12396 8432 12424
rect 8168 12384 8174 12396
rect 7561 12359 7619 12365
rect 7561 12356 7573 12359
rect 6788 12328 7328 12356
rect 7392 12328 7573 12356
rect 6788 12316 6794 12328
rect 7300 12288 7328 12328
rect 7561 12325 7573 12328
rect 7607 12356 7619 12359
rect 8294 12356 8300 12368
rect 7607 12328 8300 12356
rect 7607 12325 7619 12328
rect 7561 12319 7619 12325
rect 8294 12316 8300 12328
rect 8352 12316 8358 12368
rect 7300 12260 8340 12288
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 2314 12220 2320 12232
rect 2271 12192 2320 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 2314 12180 2320 12192
rect 2372 12220 2378 12232
rect 3326 12220 3332 12232
rect 2372 12192 3332 12220
rect 2372 12180 2378 12192
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 7098 12220 7104 12232
rect 6512 12192 7104 12220
rect 6512 12180 6518 12192
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 7650 12220 7656 12232
rect 7340 12192 7656 12220
rect 7340 12180 7346 12192
rect 7650 12180 7656 12192
rect 7708 12180 7714 12232
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 8018 12220 8024 12232
rect 7791 12192 8024 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 8202 12180 8208 12232
rect 8260 12180 8266 12232
rect 8312 12229 8340 12260
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12189 8355 12223
rect 8404 12220 8432 12396
rect 9585 12393 9597 12427
rect 9631 12424 9643 12427
rect 9674 12424 9680 12436
rect 9631 12396 9680 12424
rect 9631 12393 9643 12396
rect 9585 12387 9643 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10410 12424 10416 12436
rect 10192 12396 10416 12424
rect 10192 12384 10198 12396
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 11238 12384 11244 12436
rect 11296 12424 11302 12436
rect 11698 12424 11704 12436
rect 11296 12396 11704 12424
rect 11296 12384 11302 12396
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 15105 12427 15163 12433
rect 11940 12396 14412 12424
rect 11940 12384 11946 12396
rect 12986 12356 12992 12368
rect 9692 12328 12992 12356
rect 9692 12300 9720 12328
rect 12986 12316 12992 12328
rect 13044 12316 13050 12368
rect 14384 12300 14412 12396
rect 15105 12393 15117 12427
rect 15151 12424 15163 12427
rect 15470 12424 15476 12436
rect 15151 12396 15476 12424
rect 15151 12393 15163 12396
rect 15105 12387 15163 12393
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 16574 12424 16580 12436
rect 16356 12396 16580 12424
rect 16356 12384 16362 12396
rect 16574 12384 16580 12396
rect 16632 12384 16638 12436
rect 14645 12359 14703 12365
rect 14645 12325 14657 12359
rect 14691 12356 14703 12359
rect 15194 12356 15200 12368
rect 14691 12328 15200 12356
rect 14691 12325 14703 12328
rect 14645 12319 14703 12325
rect 15194 12316 15200 12328
rect 15252 12316 15258 12368
rect 8754 12248 8760 12300
rect 8812 12288 8818 12300
rect 8812 12260 9444 12288
rect 8812 12248 8818 12260
rect 9416 12232 9444 12260
rect 9674 12248 9680 12300
rect 9732 12248 9738 12300
rect 11422 12248 11428 12300
rect 11480 12288 11486 12300
rect 11882 12288 11888 12300
rect 11480 12260 11888 12288
rect 11480 12248 11486 12260
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 12342 12248 12348 12300
rect 12400 12288 12406 12300
rect 13357 12291 13415 12297
rect 13357 12288 13369 12291
rect 12400 12260 13369 12288
rect 12400 12248 12406 12260
rect 13357 12257 13369 12260
rect 13403 12288 13415 12291
rect 13906 12288 13912 12300
rect 13403 12260 13912 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14090 12248 14096 12300
rect 14148 12288 14154 12300
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 14148 12260 14197 12288
rect 14148 12248 14154 12260
rect 14185 12257 14197 12260
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 14366 12248 14372 12300
rect 14424 12248 14430 12300
rect 8481 12223 8539 12229
rect 8481 12220 8493 12223
rect 8404 12192 8493 12220
rect 8297 12183 8355 12189
rect 8481 12189 8493 12192
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 9398 12180 9404 12232
rect 9456 12180 9462 12232
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 4614 12112 4620 12164
rect 4672 12152 4678 12164
rect 7190 12152 7196 12164
rect 4672 12124 7196 12152
rect 4672 12112 4678 12124
rect 7190 12112 7196 12124
rect 7248 12112 7254 12164
rect 7834 12112 7840 12164
rect 7892 12152 7898 12164
rect 9508 12152 9536 12183
rect 10318 12180 10324 12232
rect 10376 12180 10382 12232
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12220 11575 12223
rect 11606 12220 11612 12232
rect 11563 12192 11612 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 11698 12180 11704 12232
rect 11756 12180 11762 12232
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 7892 12124 9536 12152
rect 7892 12112 7898 12124
rect 9508 12096 9536 12124
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10137 12155 10195 12161
rect 10137 12152 10149 12155
rect 9916 12124 10149 12152
rect 9916 12112 9922 12124
rect 10137 12121 10149 12124
rect 10183 12121 10195 12155
rect 10137 12115 10195 12121
rect 10686 12112 10692 12164
rect 10744 12112 10750 12164
rect 11808 12152 11836 12183
rect 12158 12180 12164 12232
rect 12216 12220 12222 12232
rect 12618 12220 12624 12232
rect 12216 12192 12624 12220
rect 12216 12180 12222 12192
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 12986 12180 12992 12232
rect 13044 12180 13050 12232
rect 13265 12223 13323 12229
rect 13173 12217 13231 12223
rect 13173 12183 13185 12217
rect 13219 12183 13231 12217
rect 13265 12189 13277 12223
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 13173 12177 13231 12183
rect 10980 12124 11836 12152
rect 1854 12044 1860 12096
rect 1912 12084 1918 12096
rect 2317 12087 2375 12093
rect 2317 12084 2329 12087
rect 1912 12056 2329 12084
rect 1912 12044 1918 12056
rect 2317 12053 2329 12056
rect 2363 12053 2375 12087
rect 2317 12047 2375 12053
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 6052 12056 7113 12084
rect 6052 12044 6058 12056
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 7101 12047 7159 12053
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 8202 12084 8208 12096
rect 7616 12056 8208 12084
rect 7616 12044 7622 12056
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8662 12044 8668 12096
rect 8720 12044 8726 12096
rect 9490 12044 9496 12096
rect 9548 12044 9554 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10502 12084 10508 12096
rect 9732 12056 10508 12084
rect 9732 12044 9738 12056
rect 10502 12044 10508 12056
rect 10560 12084 10566 12096
rect 10980 12084 11008 12124
rect 10560 12056 11008 12084
rect 10560 12044 10566 12056
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11422 12084 11428 12096
rect 11112 12056 11428 12084
rect 11112 12044 11118 12056
rect 11422 12044 11428 12056
rect 11480 12084 11486 12096
rect 13188 12084 13216 12177
rect 13280 12152 13308 12183
rect 13538 12180 13544 12232
rect 13596 12180 13602 12232
rect 14274 12180 14280 12232
rect 14332 12180 14338 12232
rect 14458 12180 14464 12232
rect 14516 12180 14522 12232
rect 15197 12223 15255 12229
rect 15197 12189 15209 12223
rect 15243 12220 15255 12223
rect 18046 12220 18052 12232
rect 15243 12192 18052 12220
rect 15243 12189 15255 12192
rect 15197 12183 15255 12189
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 13725 12155 13783 12161
rect 13280 12124 13492 12152
rect 13464 12096 13492 12124
rect 13725 12121 13737 12155
rect 13771 12152 13783 12155
rect 15470 12152 15476 12164
rect 13771 12124 15476 12152
rect 13771 12121 13783 12124
rect 13725 12115 13783 12121
rect 15470 12112 15476 12124
rect 15528 12112 15534 12164
rect 11480 12056 13216 12084
rect 11480 12044 11486 12056
rect 13446 12044 13452 12096
rect 13504 12044 13510 12096
rect 13906 12044 13912 12096
rect 13964 12084 13970 12096
rect 14737 12087 14795 12093
rect 14737 12084 14749 12087
rect 13964 12056 14749 12084
rect 13964 12044 13970 12056
rect 14737 12053 14749 12056
rect 14783 12053 14795 12087
rect 14737 12047 14795 12053
rect 1104 11994 18860 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 7610 11994
rect 7662 11942 7674 11994
rect 7726 11942 7738 11994
rect 7790 11942 7802 11994
rect 7854 11942 7866 11994
rect 7918 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 17610 11994
rect 17662 11942 17674 11994
rect 17726 11942 17738 11994
rect 17790 11942 17802 11994
rect 17854 11942 17866 11994
rect 17918 11942 18860 11994
rect 1104 11920 18860 11942
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 7282 11880 7288 11892
rect 4304 11852 7288 11880
rect 4304 11840 4310 11852
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 12710 11880 12716 11892
rect 7760 11852 12716 11880
rect 3786 11772 3792 11824
rect 3844 11812 3850 11824
rect 6178 11812 6184 11824
rect 3844 11784 6184 11812
rect 3844 11772 3850 11784
rect 6178 11772 6184 11784
rect 6236 11772 6242 11824
rect 7760 11812 7788 11852
rect 12710 11840 12716 11852
rect 12768 11880 12774 11892
rect 13078 11880 13084 11892
rect 12768 11852 13084 11880
rect 12768 11840 12774 11852
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 14090 11840 14096 11892
rect 14148 11880 14154 11892
rect 15378 11880 15384 11892
rect 14148 11852 15384 11880
rect 14148 11840 14154 11852
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 18690 11840 18696 11892
rect 18748 11880 18754 11892
rect 18966 11880 18972 11892
rect 18748 11852 18972 11880
rect 18748 11840 18754 11852
rect 18966 11840 18972 11852
rect 19024 11840 19030 11892
rect 7576 11784 7788 11812
rect 842 11704 848 11756
rect 900 11744 906 11756
rect 1489 11747 1547 11753
rect 1489 11744 1501 11747
rect 900 11716 1501 11744
rect 900 11704 906 11716
rect 1489 11713 1501 11716
rect 1535 11713 1547 11747
rect 1489 11707 1547 11713
rect 3881 11747 3939 11753
rect 3881 11713 3893 11747
rect 3927 11713 3939 11747
rect 3881 11707 3939 11713
rect 3973 11747 4031 11753
rect 3973 11713 3985 11747
rect 4019 11744 4031 11747
rect 5810 11744 5816 11756
rect 4019 11716 5816 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 3896 11676 3924 11707
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 6454 11744 6460 11756
rect 5960 11716 6460 11744
rect 5960 11704 5966 11716
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 4062 11676 4068 11688
rect 3896 11648 4068 11676
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 7208 11676 7236 11707
rect 7282 11704 7288 11756
rect 7340 11704 7346 11756
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11744 7527 11747
rect 7576 11744 7604 11784
rect 7834 11772 7840 11824
rect 7892 11812 7898 11824
rect 9582 11812 9588 11824
rect 7892 11784 9588 11812
rect 7892 11772 7898 11784
rect 9582 11772 9588 11784
rect 9640 11812 9646 11824
rect 9640 11784 11836 11812
rect 9640 11772 9646 11784
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 7515 11716 7604 11744
rect 7668 11716 10333 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 7558 11676 7564 11688
rect 7208 11648 7564 11676
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 1673 11611 1731 11617
rect 1673 11577 1685 11611
rect 1719 11608 1731 11611
rect 2958 11608 2964 11620
rect 1719 11580 2964 11608
rect 1719 11577 1731 11580
rect 1673 11571 1731 11577
rect 2958 11568 2964 11580
rect 3016 11608 3022 11620
rect 7668 11608 7696 11716
rect 10321 11713 10333 11716
rect 10367 11744 10379 11747
rect 10594 11744 10600 11756
rect 10367 11716 10600 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 7742 11636 7748 11688
rect 7800 11676 7806 11688
rect 8478 11676 8484 11688
rect 7800 11648 8484 11676
rect 7800 11636 7806 11648
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 10226 11636 10232 11688
rect 10284 11636 10290 11688
rect 11808 11676 11836 11784
rect 11974 11772 11980 11824
rect 12032 11812 12038 11824
rect 12032 11784 12434 11812
rect 12032 11772 12038 11784
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 11940 11716 12173 11744
rect 11940 11704 11946 11716
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12406 11744 12434 11784
rect 13170 11772 13176 11824
rect 13228 11812 13234 11824
rect 13630 11812 13636 11824
rect 13228 11784 13636 11812
rect 13228 11772 13234 11784
rect 13630 11772 13636 11784
rect 13688 11772 13694 11824
rect 14274 11772 14280 11824
rect 14332 11772 14338 11824
rect 14550 11812 14556 11824
rect 14476 11784 14556 11812
rect 14182 11744 14188 11756
rect 12406 11716 14188 11744
rect 12161 11707 12219 11713
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 14476 11753 14504 11784
rect 14550 11772 14556 11784
rect 14608 11812 14614 11824
rect 15102 11812 15108 11824
rect 14608 11784 15108 11812
rect 14608 11772 14614 11784
rect 15102 11772 15108 11784
rect 15160 11772 15166 11824
rect 14461 11747 14519 11753
rect 14461 11713 14473 11747
rect 14507 11713 14519 11747
rect 14461 11707 14519 11713
rect 14645 11747 14703 11753
rect 14645 11713 14657 11747
rect 14691 11713 14703 11747
rect 14645 11707 14703 11713
rect 14660 11676 14688 11707
rect 15378 11704 15384 11756
rect 15436 11744 15442 11756
rect 17773 11747 17831 11753
rect 17773 11744 17785 11747
rect 15436 11716 17785 11744
rect 15436 11704 15442 11716
rect 17773 11713 17785 11716
rect 17819 11713 17831 11747
rect 17773 11707 17831 11713
rect 18233 11747 18291 11753
rect 18233 11713 18245 11747
rect 18279 11744 18291 11747
rect 18690 11744 18696 11756
rect 18279 11716 18696 11744
rect 18279 11713 18291 11716
rect 18233 11707 18291 11713
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 15838 11676 15844 11688
rect 11808 11648 14596 11676
rect 14660 11648 15844 11676
rect 3016 11580 7696 11608
rect 3016 11568 3022 11580
rect 8202 11568 8208 11620
rect 8260 11608 8266 11620
rect 11606 11608 11612 11620
rect 8260 11580 11612 11608
rect 8260 11568 8266 11580
rect 11606 11568 11612 11580
rect 11664 11608 11670 11620
rect 12158 11608 12164 11620
rect 11664 11580 12164 11608
rect 11664 11568 11670 11580
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 14568 11608 14596 11648
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 17310 11636 17316 11688
rect 17368 11676 17374 11688
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 17368 11648 17509 11676
rect 17368 11636 17374 11648
rect 17497 11645 17509 11648
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 17589 11679 17647 11685
rect 17589 11645 17601 11679
rect 17635 11645 17647 11679
rect 17589 11639 17647 11645
rect 17681 11679 17739 11685
rect 17681 11645 17693 11679
rect 17727 11676 17739 11679
rect 18138 11676 18144 11688
rect 17727 11648 18144 11676
rect 17727 11645 17739 11648
rect 17681 11639 17739 11645
rect 14826 11608 14832 11620
rect 14568 11580 14832 11608
rect 14826 11568 14832 11580
rect 14884 11568 14890 11620
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 17604 11608 17632 11639
rect 18138 11636 18144 11648
rect 18196 11636 18202 11688
rect 15068 11580 17632 11608
rect 17957 11611 18015 11617
rect 15068 11568 15074 11580
rect 17957 11577 17969 11611
rect 18003 11608 18015 11611
rect 18598 11608 18604 11620
rect 18003 11580 18604 11608
rect 18003 11577 18015 11580
rect 17957 11571 18015 11577
rect 18598 11568 18604 11580
rect 18656 11568 18662 11620
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 2314 11540 2320 11552
rect 1544 11512 2320 11540
rect 1544 11500 1550 11512
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 3970 11500 3976 11552
rect 4028 11500 4034 11552
rect 5810 11500 5816 11552
rect 5868 11540 5874 11552
rect 6546 11540 6552 11552
rect 5868 11512 6552 11540
rect 5868 11500 5874 11512
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7558 11540 7564 11552
rect 7156 11512 7564 11540
rect 7156 11500 7162 11512
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 7650 11500 7656 11552
rect 7708 11500 7714 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 10045 11543 10103 11549
rect 10045 11540 10057 11543
rect 8904 11512 10057 11540
rect 8904 11500 8910 11512
rect 10045 11509 10057 11512
rect 10091 11540 10103 11543
rect 10962 11540 10968 11552
rect 10091 11512 10968 11540
rect 10091 11509 10103 11512
rect 10045 11503 10103 11509
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11514 11500 11520 11552
rect 11572 11540 11578 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11572 11512 11805 11540
rect 11572 11500 11578 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 12618 11540 12624 11552
rect 12124 11512 12624 11540
rect 12124 11500 12130 11512
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13262 11540 13268 11552
rect 13044 11512 13268 11540
rect 13044 11500 13050 11512
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 16114 11540 16120 11552
rect 14424 11512 16120 11540
rect 14424 11500 14430 11512
rect 16114 11500 16120 11512
rect 16172 11500 16178 11552
rect 18414 11500 18420 11552
rect 18472 11500 18478 11552
rect 1104 11450 18860 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 11950 11450
rect 12002 11398 12014 11450
rect 12066 11398 12078 11450
rect 12130 11398 12142 11450
rect 12194 11398 12206 11450
rect 12258 11398 16950 11450
rect 17002 11398 17014 11450
rect 17066 11398 17078 11450
rect 17130 11398 17142 11450
rect 17194 11398 17206 11450
rect 17258 11398 18860 11450
rect 1104 11376 18860 11398
rect 3326 11296 3332 11348
rect 3384 11336 3390 11348
rect 3384 11308 5856 11336
rect 3384 11296 3390 11308
rect 1486 11228 1492 11280
rect 1544 11268 1550 11280
rect 1670 11268 1676 11280
rect 1544 11240 1676 11268
rect 1544 11228 1550 11240
rect 1670 11228 1676 11240
rect 1728 11228 1734 11280
rect 3786 11268 3792 11280
rect 2148 11240 3792 11268
rect 2148 11209 2176 11240
rect 3786 11228 3792 11240
rect 3844 11228 3850 11280
rect 5534 11268 5540 11280
rect 4172 11240 5540 11268
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11169 2191 11203
rect 2133 11163 2191 11169
rect 1670 11092 1676 11144
rect 1728 11132 1734 11144
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 1728 11104 2329 11132
rect 1728 11092 1734 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11101 2559 11135
rect 2501 11095 2559 11101
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11132 2651 11135
rect 4172 11132 4200 11240
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 4706 11200 4712 11212
rect 4448 11172 4712 11200
rect 4448 11144 4476 11172
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5828 11200 5856 11308
rect 5902 11296 5908 11348
rect 5960 11296 5966 11348
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 7282 11336 7288 11348
rect 6512 11308 7288 11336
rect 6512 11296 6518 11308
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 9030 11336 9036 11348
rect 8904 11308 9036 11336
rect 8904 11296 8910 11308
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 9214 11296 9220 11348
rect 9272 11336 9278 11348
rect 9272 11308 14964 11336
rect 9272 11296 9278 11308
rect 7650 11228 7656 11280
rect 7708 11268 7714 11280
rect 14550 11268 14556 11280
rect 7708 11240 14320 11268
rect 7708 11228 7714 11240
rect 5828 11172 6684 11200
rect 2639 11104 4200 11132
rect 2639 11101 2651 11104
rect 2593 11095 2651 11101
rect 2516 11064 2544 11095
rect 4430 11092 4436 11144
rect 4488 11092 4494 11144
rect 4798 11092 4804 11144
rect 4856 11092 4862 11144
rect 5077 11135 5135 11141
rect 5077 11132 5089 11135
rect 5000 11104 5089 11132
rect 4338 11064 4344 11076
rect 2516 11036 4344 11064
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 5000 10996 5028 11104
rect 5077 11101 5089 11104
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5718 11092 5724 11144
rect 5776 11132 5782 11144
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5776 11104 5917 11132
rect 5776 11092 5782 11104
rect 5905 11101 5917 11104
rect 5951 11101 5963 11135
rect 5905 11095 5963 11101
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11132 6055 11135
rect 6656 11132 6684 11172
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 7524 11172 12480 11200
rect 7524 11160 7530 11172
rect 9858 11132 9864 11144
rect 6043 11104 6132 11132
rect 6656 11104 9864 11132
rect 6043 11101 6055 11104
rect 5997 11095 6055 11101
rect 5350 11024 5356 11076
rect 5408 11024 5414 11076
rect 6104 11008 6132 11104
rect 9858 11092 9864 11104
rect 9916 11092 9922 11144
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11514 11132 11520 11144
rect 11112 11104 11520 11132
rect 11112 11092 11118 11104
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 12250 11132 12256 11144
rect 11848 11104 12256 11132
rect 11848 11092 11854 11104
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 12342 11092 12348 11144
rect 12400 11092 12406 11144
rect 12452 11132 12480 11172
rect 12526 11160 12532 11212
rect 12584 11160 12590 11212
rect 14292 11209 14320 11240
rect 14476 11240 14556 11268
rect 14476 11209 14504 11240
rect 14550 11228 14556 11240
rect 14608 11228 14614 11280
rect 14936 11268 14964 11308
rect 15286 11296 15292 11348
rect 15344 11296 15350 11348
rect 16206 11336 16212 11348
rect 15396 11308 16212 11336
rect 15396 11268 15424 11308
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 14936 11240 15424 11268
rect 14093 11203 14151 11209
rect 14093 11169 14105 11203
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 14108 11132 14136 11163
rect 14826 11160 14832 11212
rect 14884 11160 14890 11212
rect 14936 11209 14964 11240
rect 15562 11228 15568 11280
rect 15620 11268 15626 11280
rect 16025 11271 16083 11277
rect 16025 11268 16037 11271
rect 15620 11240 16037 11268
rect 15620 11228 15626 11240
rect 16025 11237 16037 11240
rect 16071 11237 16083 11271
rect 16025 11231 16083 11237
rect 14921 11203 14979 11209
rect 14921 11169 14933 11203
rect 14967 11169 14979 11203
rect 14921 11163 14979 11169
rect 15010 11160 15016 11212
rect 15068 11160 15074 11212
rect 15105 11203 15163 11209
rect 15105 11169 15117 11203
rect 15151 11200 15163 11203
rect 15930 11200 15936 11212
rect 15151 11172 15936 11200
rect 15151 11169 15163 11172
rect 15105 11163 15163 11169
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 12452 11104 14136 11132
rect 14182 11092 14188 11144
rect 14240 11132 14246 11144
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 14240 11104 14381 11132
rect 14240 11092 14246 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11101 14611 11135
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 14553 11095 14611 11101
rect 15120 11104 16221 11132
rect 10870 11024 10876 11076
rect 10928 11064 10934 11076
rect 14568 11064 14596 11095
rect 10928 11036 14596 11064
rect 10928 11024 10934 11036
rect 14642 11024 14648 11076
rect 14700 11064 14706 11076
rect 14826 11064 14832 11076
rect 14700 11036 14832 11064
rect 14700 11024 14706 11036
rect 14826 11024 14832 11036
rect 14884 11064 14890 11076
rect 15120 11064 15148 11104
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 15933 11067 15991 11073
rect 15933 11064 15945 11067
rect 14884 11036 15148 11064
rect 15212 11036 15945 11064
rect 14884 11024 14890 11036
rect 4028 10968 5028 10996
rect 4028 10956 4034 10968
rect 6086 10956 6092 11008
rect 6144 10956 6150 11008
rect 6273 10999 6331 11005
rect 6273 10965 6285 10999
rect 6319 10996 6331 10999
rect 6454 10996 6460 11008
rect 6319 10968 6460 10996
rect 6319 10965 6331 10968
rect 6273 10959 6331 10965
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 12529 10999 12587 11005
rect 12529 10965 12541 10999
rect 12575 10996 12587 10999
rect 12618 10996 12624 11008
rect 12575 10968 12624 10996
rect 12575 10965 12587 10968
rect 12529 10959 12587 10965
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 13262 10956 13268 11008
rect 13320 10996 13326 11008
rect 14090 10996 14096 11008
rect 13320 10968 14096 10996
rect 13320 10956 13326 10968
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 14458 10956 14464 11008
rect 14516 10996 14522 11008
rect 15212 10996 15240 11036
rect 15933 11033 15945 11036
rect 15979 11033 15991 11067
rect 15933 11027 15991 11033
rect 16114 11024 16120 11076
rect 16172 11024 16178 11076
rect 14516 10968 15240 10996
rect 14516 10956 14522 10968
rect 1104 10906 18860 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 17610 10906
rect 17662 10854 17674 10906
rect 17726 10854 17738 10906
rect 17790 10854 17802 10906
rect 17854 10854 17866 10906
rect 17918 10854 18860 10906
rect 1104 10832 18860 10854
rect 3970 10752 3976 10804
rect 4028 10752 4034 10804
rect 4065 10795 4123 10801
rect 4065 10761 4077 10795
rect 4111 10792 4123 10795
rect 4154 10792 4160 10804
rect 4111 10764 4160 10792
rect 4111 10761 4123 10764
rect 4065 10755 4123 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4522 10792 4528 10804
rect 4356 10764 4528 10792
rect 1489 10727 1547 10733
rect 1489 10693 1501 10727
rect 1535 10724 1547 10727
rect 1578 10724 1584 10736
rect 1535 10696 1584 10724
rect 1535 10693 1547 10696
rect 1489 10687 1547 10693
rect 1578 10684 1584 10696
rect 1636 10684 1642 10736
rect 3786 10684 3792 10736
rect 3844 10684 3850 10736
rect 3988 10724 4016 10752
rect 4356 10733 4384 10764
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 4709 10795 4767 10801
rect 4709 10761 4721 10795
rect 4755 10792 4767 10795
rect 4755 10764 4936 10792
rect 4755 10761 4767 10764
rect 4709 10755 4767 10761
rect 4341 10727 4399 10733
rect 3896 10696 4292 10724
rect 1670 10616 1676 10668
rect 1728 10616 1734 10668
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 1854 10656 1860 10668
rect 1811 10628 1860 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 1854 10616 1860 10628
rect 1912 10616 1918 10668
rect 1946 10616 1952 10668
rect 2004 10616 2010 10668
rect 3510 10656 3516 10668
rect 2746 10628 3516 10656
rect 1872 10520 1900 10616
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2746 10588 2774 10628
rect 3510 10616 3516 10628
rect 3568 10656 3574 10668
rect 3896 10656 3924 10696
rect 3568 10628 3924 10656
rect 3568 10616 3574 10628
rect 3970 10616 3976 10668
rect 4028 10616 4034 10668
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4264 10656 4292 10696
rect 4341 10693 4353 10727
rect 4387 10693 4399 10727
rect 4341 10687 4399 10693
rect 4614 10684 4620 10736
rect 4672 10724 4678 10736
rect 4801 10727 4859 10733
rect 4801 10724 4813 10727
rect 4672 10696 4813 10724
rect 4672 10684 4678 10696
rect 4801 10693 4813 10696
rect 4847 10693 4859 10727
rect 4908 10724 4936 10764
rect 4982 10752 4988 10804
rect 5040 10752 5046 10804
rect 5350 10752 5356 10804
rect 5408 10792 5414 10804
rect 9030 10792 9036 10804
rect 5408 10764 9036 10792
rect 5408 10752 5414 10764
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 15102 10792 15108 10804
rect 9180 10764 15108 10792
rect 9180 10752 9186 10764
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 15194 10724 15200 10736
rect 4908 10696 15200 10724
rect 4801 10687 4859 10693
rect 15194 10684 15200 10696
rect 15252 10684 15258 10736
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4264 10628 4445 10656
rect 4157 10619 4215 10625
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10656 4583 10659
rect 5074 10656 5080 10668
rect 4571 10628 5080 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 2271 10560 2774 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 3418 10588 3424 10600
rect 3108 10560 3424 10588
rect 3108 10548 3114 10560
rect 3418 10548 3424 10560
rect 3476 10588 3482 10600
rect 4080 10588 4108 10619
rect 3476 10560 4108 10588
rect 4172 10588 4200 10619
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 8754 10656 8760 10668
rect 5307 10628 8760 10656
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 12526 10656 12532 10668
rect 12308 10628 12532 10656
rect 12308 10616 12314 10628
rect 12526 10616 12532 10628
rect 12584 10656 12590 10668
rect 13630 10656 13636 10668
rect 12584 10628 13636 10656
rect 12584 10616 12590 10628
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10625 13783 10659
rect 13725 10619 13783 10625
rect 4706 10588 4712 10600
rect 4172 10560 4712 10588
rect 3476 10548 3482 10560
rect 4172 10520 4200 10560
rect 4706 10548 4712 10560
rect 4764 10588 4770 10600
rect 9950 10588 9956 10600
rect 4764 10560 9956 10588
rect 4764 10548 4770 10560
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 13262 10548 13268 10600
rect 13320 10588 13326 10600
rect 13740 10588 13768 10619
rect 13814 10616 13820 10668
rect 13872 10616 13878 10668
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10656 14151 10659
rect 14182 10656 14188 10668
rect 14139 10628 14188 10656
rect 14139 10625 14151 10628
rect 14093 10619 14151 10625
rect 14182 10616 14188 10628
rect 14240 10616 14246 10668
rect 15010 10616 15016 10668
rect 15068 10656 15074 10668
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 15068 10628 18245 10656
rect 15068 10616 15074 10628
rect 18233 10625 18245 10628
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 13320 10560 13768 10588
rect 14277 10591 14335 10597
rect 13320 10548 13326 10560
rect 14277 10557 14289 10591
rect 14323 10588 14335 10591
rect 14642 10588 14648 10600
rect 14323 10560 14648 10588
rect 14323 10557 14335 10560
rect 14277 10551 14335 10557
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15378 10588 15384 10600
rect 14976 10560 15384 10588
rect 14976 10548 14982 10560
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 1872 10492 4200 10520
rect 4522 10480 4528 10532
rect 4580 10520 4586 10532
rect 4890 10520 4896 10532
rect 4580 10492 4896 10520
rect 4580 10480 4586 10492
rect 4890 10480 4896 10492
rect 4948 10480 4954 10532
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 12618 10520 12624 10532
rect 5408 10492 12624 10520
rect 5408 10480 5414 10492
rect 12618 10480 12624 10492
rect 12676 10520 12682 10532
rect 17954 10520 17960 10532
rect 12676 10492 17960 10520
rect 12676 10480 12682 10492
rect 17954 10480 17960 10492
rect 18012 10480 18018 10532
rect 1486 10412 1492 10464
rect 1544 10412 1550 10464
rect 4985 10455 5043 10461
rect 4985 10421 4997 10455
rect 5031 10452 5043 10455
rect 11790 10452 11796 10464
rect 5031 10424 11796 10452
rect 5031 10421 5043 10424
rect 4985 10415 5043 10421
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 13998 10412 14004 10464
rect 14056 10452 14062 10464
rect 17770 10452 17776 10464
rect 14056 10424 17776 10452
rect 14056 10412 14062 10424
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 18414 10412 18420 10464
rect 18472 10412 18478 10464
rect 1104 10362 18860 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 11950 10362
rect 12002 10310 12014 10362
rect 12066 10310 12078 10362
rect 12130 10310 12142 10362
rect 12194 10310 12206 10362
rect 12258 10310 16950 10362
rect 17002 10310 17014 10362
rect 17066 10310 17078 10362
rect 17130 10310 17142 10362
rect 17194 10310 17206 10362
rect 17258 10310 18860 10362
rect 1104 10288 18860 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 17589 10251 17647 10257
rect 17589 10248 17601 10251
rect 1544 10220 4844 10248
rect 1544 10208 1550 10220
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 1719 10084 4752 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 842 10004 848 10056
rect 900 10044 906 10056
rect 1489 10047 1547 10053
rect 1489 10044 1501 10047
rect 900 10016 1501 10044
rect 900 10004 906 10016
rect 1489 10013 1501 10016
rect 1535 10013 1547 10047
rect 1489 10007 1547 10013
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 1857 10047 1915 10053
rect 1857 10044 1869 10047
rect 1820 10016 1869 10044
rect 1820 10004 1826 10016
rect 1857 10013 1869 10016
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10013 2099 10047
rect 2041 10007 2099 10013
rect 1578 9936 1584 9988
rect 1636 9976 1642 9988
rect 2056 9976 2084 10007
rect 1636 9948 2084 9976
rect 1636 9936 1642 9948
rect 1949 9911 2007 9917
rect 1949 9877 1961 9911
rect 1995 9908 2007 9911
rect 3694 9908 3700 9920
rect 1995 9880 3700 9908
rect 1995 9877 2007 9880
rect 1949 9871 2007 9877
rect 3694 9868 3700 9880
rect 3752 9908 3758 9920
rect 4062 9908 4068 9920
rect 3752 9880 4068 9908
rect 3752 9868 3758 9880
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4724 9908 4752 10084
rect 4816 9976 4844 10220
rect 4908 10220 17601 10248
rect 4908 10053 4936 10220
rect 17589 10217 17601 10220
rect 17635 10217 17647 10251
rect 17589 10211 17647 10217
rect 17770 10208 17776 10260
rect 17828 10208 17834 10260
rect 4982 10140 4988 10192
rect 5040 10140 5046 10192
rect 5074 10140 5080 10192
rect 5132 10140 5138 10192
rect 11146 10180 11152 10192
rect 10704 10152 11152 10180
rect 5000 10112 5028 10140
rect 7558 10112 7564 10124
rect 5000 10084 7564 10112
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 10704 10121 10732 10152
rect 11146 10140 11152 10152
rect 11204 10140 11210 10192
rect 14918 10180 14924 10192
rect 11440 10152 14924 10180
rect 10689 10115 10747 10121
rect 10689 10081 10701 10115
rect 10735 10081 10747 10115
rect 10689 10075 10747 10081
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 5040 10016 10548 10044
rect 5040 10004 5046 10016
rect 9766 9976 9772 9988
rect 4816 9948 9772 9976
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 10520 9976 10548 10016
rect 10594 10004 10600 10056
rect 10652 10004 10658 10056
rect 11440 10053 11468 10152
rect 14918 10140 14924 10152
rect 14976 10140 14982 10192
rect 15013 10183 15071 10189
rect 15013 10149 15025 10183
rect 15059 10180 15071 10183
rect 15378 10180 15384 10192
rect 15059 10152 15384 10180
rect 15059 10149 15071 10152
rect 15013 10143 15071 10149
rect 15378 10140 15384 10152
rect 15436 10140 15442 10192
rect 16574 10140 16580 10192
rect 16632 10180 16638 10192
rect 17954 10180 17960 10192
rect 16632 10152 16988 10180
rect 16632 10140 16638 10152
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10112 11851 10115
rect 12618 10112 12624 10124
rect 11839 10084 12624 10112
rect 11839 10081 11851 10084
rect 11793 10075 11851 10081
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 13630 10072 13636 10124
rect 13688 10112 13694 10124
rect 15396 10112 15424 10140
rect 16850 10112 16856 10124
rect 13688 10084 14872 10112
rect 15396 10084 16856 10112
rect 13688 10072 13694 10084
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 11072 10016 11437 10044
rect 11072 9976 11100 10016
rect 11425 10013 11437 10016
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10044 11759 10047
rect 11882 10044 11888 10056
rect 11747 10016 11888 10044
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 11882 10004 11888 10016
rect 11940 10044 11946 10056
rect 13998 10044 14004 10056
rect 11940 10016 14004 10044
rect 11940 10004 11946 10016
rect 13998 10004 14004 10016
rect 14056 10044 14062 10056
rect 14645 10047 14703 10053
rect 14645 10044 14657 10047
rect 14056 10016 14657 10044
rect 14056 10004 14062 10016
rect 14645 10013 14657 10016
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 10520 9948 11100 9976
rect 11330 9936 11336 9988
rect 11388 9976 11394 9988
rect 13814 9976 13820 9988
rect 11388 9948 13820 9976
rect 11388 9936 11394 9948
rect 13814 9936 13820 9948
rect 13872 9976 13878 9988
rect 14737 9979 14795 9985
rect 14737 9976 14749 9979
rect 13872 9948 14749 9976
rect 13872 9936 13878 9948
rect 14737 9945 14749 9948
rect 14783 9945 14795 9979
rect 14737 9939 14795 9945
rect 8202 9908 8208 9920
rect 4724 9880 8208 9908
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 10962 9868 10968 9920
rect 11020 9868 11026 9920
rect 14274 9868 14280 9920
rect 14332 9908 14338 9920
rect 14844 9917 14872 10084
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 15102 10004 15108 10056
rect 15160 10004 15166 10056
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 16960 10053 16988 10152
rect 17420 10152 17960 10180
rect 17420 10121 17448 10152
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 17862 10072 17868 10124
rect 17920 10072 17926 10124
rect 16577 10047 16635 10053
rect 16577 10044 16589 10047
rect 15252 10016 16589 10044
rect 15252 10004 15258 10016
rect 16577 10013 16589 10016
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10013 17831 10047
rect 17773 10007 17831 10013
rect 15378 9936 15384 9988
rect 15436 9936 15442 9988
rect 16390 9936 16396 9988
rect 16448 9936 16454 9988
rect 17034 9936 17040 9988
rect 17092 9976 17098 9988
rect 17788 9976 17816 10007
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 17092 9948 17816 9976
rect 17092 9936 17098 9948
rect 14461 9911 14519 9917
rect 14461 9908 14473 9911
rect 14332 9880 14473 9908
rect 14332 9868 14338 9880
rect 14461 9877 14473 9880
rect 14507 9877 14519 9911
rect 14461 9871 14519 9877
rect 14829 9911 14887 9917
rect 14829 9877 14841 9911
rect 14875 9908 14887 9911
rect 18414 9908 18420 9920
rect 14875 9880 18420 9908
rect 14875 9877 14887 9880
rect 14829 9871 14887 9877
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 1104 9818 18860 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 17610 9818
rect 17662 9766 17674 9818
rect 17726 9766 17738 9818
rect 17790 9766 17802 9818
rect 17854 9766 17866 9818
rect 17918 9766 18860 9818
rect 1104 9744 18860 9766
rect 1581 9707 1639 9713
rect 1581 9673 1593 9707
rect 1627 9673 1639 9707
rect 3142 9704 3148 9716
rect 1581 9667 1639 9673
rect 2976 9676 3148 9704
rect 1596 9636 1624 9667
rect 2976 9636 3004 9676
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 5350 9664 5356 9716
rect 5408 9713 5414 9716
rect 5408 9707 5427 9713
rect 5415 9673 5427 9707
rect 5408 9667 5427 9673
rect 5408 9664 5414 9667
rect 7282 9664 7288 9716
rect 7340 9704 7346 9716
rect 8294 9704 8300 9716
rect 7340 9676 8300 9704
rect 7340 9664 7346 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 11882 9704 11888 9716
rect 10008 9676 11888 9704
rect 10008 9664 10014 9676
rect 11882 9664 11888 9676
rect 11940 9664 11946 9716
rect 13722 9664 13728 9716
rect 13780 9704 13786 9716
rect 15378 9704 15384 9716
rect 13780 9676 15384 9704
rect 13780 9664 13786 9676
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 16022 9664 16028 9716
rect 16080 9704 16086 9716
rect 16080 9676 16160 9704
rect 16080 9664 16086 9676
rect 16132 9674 16160 9676
rect 1596 9608 3004 9636
rect 3050 9596 3056 9648
rect 3108 9636 3114 9648
rect 3237 9639 3295 9645
rect 3237 9636 3249 9639
rect 3108 9608 3249 9636
rect 3108 9596 3114 9608
rect 3237 9605 3249 9608
rect 3283 9605 3295 9639
rect 3237 9599 3295 9605
rect 5169 9639 5227 9645
rect 5169 9605 5181 9639
rect 5215 9636 5227 9639
rect 5258 9636 5264 9648
rect 5215 9608 5264 9636
rect 5215 9605 5227 9608
rect 5169 9599 5227 9605
rect 5258 9596 5264 9608
rect 5316 9596 5322 9648
rect 10042 9636 10048 9648
rect 5460 9608 10048 9636
rect 842 9528 848 9580
rect 900 9568 906 9580
rect 1397 9571 1455 9577
rect 1397 9568 1409 9571
rect 900 9540 1409 9568
rect 900 9528 906 9540
rect 1397 9537 1409 9540
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2222 9568 2228 9580
rect 2087 9540 2228 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 2866 9568 2872 9580
rect 2455 9540 2872 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2332 9432 2360 9531
rect 2866 9528 2872 9540
rect 2924 9528 2930 9580
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 2976 9500 3004 9531
rect 3142 9528 3148 9580
rect 3200 9528 3206 9580
rect 3326 9528 3332 9580
rect 3384 9528 3390 9580
rect 4522 9500 4528 9512
rect 2976 9472 4528 9500
rect 4522 9460 4528 9472
rect 4580 9500 4586 9512
rect 5460 9500 5488 9608
rect 10042 9596 10048 9608
rect 10100 9596 10106 9648
rect 16132 9646 16436 9674
rect 16574 9664 16580 9716
rect 16632 9664 16638 9716
rect 16758 9664 16764 9716
rect 16816 9664 16822 9716
rect 5994 9528 6000 9580
rect 6052 9528 6058 9580
rect 6086 9528 6092 9580
rect 6144 9568 6150 9580
rect 6638 9568 6644 9580
rect 6144 9540 6644 9568
rect 6144 9528 6150 9540
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 9674 9568 9680 9580
rect 6972 9540 9680 9568
rect 6972 9528 6978 9540
rect 9674 9528 9680 9540
rect 9732 9568 9738 9580
rect 10778 9568 10784 9580
rect 9732 9540 10784 9568
rect 9732 9528 9738 9540
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 15378 9568 15384 9580
rect 15252 9540 15384 9568
rect 15252 9528 15258 9540
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 15746 9528 15752 9580
rect 15804 9568 15810 9580
rect 16197 9569 16255 9575
rect 15804 9566 16160 9568
rect 16197 9566 16209 9569
rect 15804 9540 16209 9566
rect 15804 9528 15810 9540
rect 16132 9538 16209 9540
rect 16197 9535 16209 9538
rect 16243 9535 16255 9569
rect 16408 9568 16436 9646
rect 16592 9636 16620 9664
rect 16197 9529 16255 9535
rect 16316 9540 16436 9568
rect 16500 9608 16620 9636
rect 16776 9636 16804 9664
rect 18417 9639 18475 9645
rect 18417 9636 18429 9639
rect 16776 9608 18429 9636
rect 4580 9472 5488 9500
rect 4580 9460 4586 9472
rect 5718 9460 5724 9512
rect 5776 9460 5782 9512
rect 5810 9460 5816 9512
rect 5868 9460 5874 9512
rect 5902 9460 5908 9512
rect 5960 9460 5966 9512
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 6512 9472 8984 9500
rect 6512 9460 6518 9472
rect 3513 9435 3571 9441
rect 2332 9404 2774 9432
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 2133 9367 2191 9373
rect 2133 9364 2145 9367
rect 1912 9336 2145 9364
rect 1912 9324 1918 9336
rect 2133 9333 2145 9336
rect 2179 9333 2191 9367
rect 2133 9327 2191 9333
rect 2590 9324 2596 9376
rect 2648 9324 2654 9376
rect 2746 9364 2774 9404
rect 3513 9401 3525 9435
rect 3559 9432 3571 9435
rect 3602 9432 3608 9444
rect 3559 9404 3608 9432
rect 3559 9401 3571 9404
rect 3513 9395 3571 9401
rect 3602 9392 3608 9404
rect 3660 9392 3666 9444
rect 3970 9392 3976 9444
rect 4028 9432 4034 9444
rect 5537 9435 5595 9441
rect 4028 9404 5396 9432
rect 4028 9392 4034 9404
rect 5074 9364 5080 9376
rect 2746 9336 5080 9364
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5368 9373 5396 9404
rect 5537 9401 5549 9435
rect 5583 9432 5595 9435
rect 5626 9432 5632 9444
rect 5583 9404 5632 9432
rect 5583 9401 5595 9404
rect 5537 9395 5595 9401
rect 5626 9392 5632 9404
rect 5684 9392 5690 9444
rect 6638 9432 6644 9444
rect 5736 9404 6644 9432
rect 5353 9367 5411 9373
rect 5353 9333 5365 9367
rect 5399 9364 5411 9367
rect 5736 9364 5764 9404
rect 6638 9392 6644 9404
rect 6696 9392 6702 9444
rect 8956 9432 8984 9472
rect 9030 9460 9036 9512
rect 9088 9500 9094 9512
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 9088 9472 16037 9500
rect 9088 9460 9094 9472
rect 16025 9469 16037 9472
rect 16071 9500 16083 9503
rect 16316 9500 16344 9540
rect 16500 9500 16528 9608
rect 18417 9605 18429 9608
rect 18463 9605 18475 9639
rect 18417 9599 18475 9605
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16632 9540 16681 9568
rect 16632 9528 16638 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 16071 9472 16344 9500
rect 16408 9472 16528 9500
rect 16868 9500 16896 9531
rect 16942 9528 16948 9580
rect 17000 9568 17006 9580
rect 17957 9571 18015 9577
rect 17957 9568 17969 9571
rect 17000 9540 17969 9568
rect 17000 9528 17006 9540
rect 17957 9537 17969 9540
rect 18003 9537 18015 9571
rect 17957 9531 18015 9537
rect 18322 9528 18328 9580
rect 18380 9528 18386 9580
rect 17126 9500 17132 9512
rect 16868 9472 17132 9500
rect 16071 9469 16083 9472
rect 16025 9463 16083 9469
rect 10410 9432 10416 9444
rect 8956 9404 10416 9432
rect 10410 9392 10416 9404
rect 10468 9432 10474 9444
rect 15010 9432 15016 9444
rect 10468 9404 15016 9432
rect 10468 9392 10474 9404
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 5399 9336 5764 9364
rect 6181 9367 6239 9373
rect 5399 9333 5411 9336
rect 5353 9327 5411 9333
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 15930 9364 15936 9376
rect 6227 9336 15936 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16408 9373 16436 9472
rect 17126 9460 17132 9472
rect 17184 9500 17190 9512
rect 17862 9500 17868 9512
rect 17184 9472 17868 9500
rect 17184 9460 17190 9472
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 18230 9460 18236 9512
rect 18288 9460 18294 9512
rect 18049 9435 18107 9441
rect 18049 9401 18061 9435
rect 18095 9432 18107 9435
rect 18414 9432 18420 9444
rect 18095 9404 18420 9432
rect 18095 9401 18107 9404
rect 18049 9395 18107 9401
rect 18414 9392 18420 9404
rect 18472 9392 18478 9444
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 16356 9336 16405 9364
rect 16356 9324 16362 9336
rect 16393 9333 16405 9336
rect 16439 9333 16451 9367
rect 16393 9327 16451 9333
rect 16761 9367 16819 9373
rect 16761 9333 16773 9367
rect 16807 9364 16819 9367
rect 17586 9364 17592 9376
rect 16807 9336 17592 9364
rect 16807 9333 16819 9336
rect 16761 9327 16819 9333
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 1104 9274 18860 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 11950 9274
rect 12002 9222 12014 9274
rect 12066 9222 12078 9274
rect 12130 9222 12142 9274
rect 12194 9222 12206 9274
rect 12258 9222 16950 9274
rect 17002 9222 17014 9274
rect 17066 9222 17078 9274
rect 17130 9222 17142 9274
rect 17194 9222 17206 9274
rect 17258 9222 18860 9274
rect 1104 9200 18860 9222
rect 2133 9163 2191 9169
rect 2133 9129 2145 9163
rect 2179 9160 2191 9163
rect 5534 9160 5540 9172
rect 2179 9132 5540 9160
rect 2179 9129 2191 9132
rect 2133 9123 2191 9129
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 13078 9160 13084 9172
rect 5868 9132 13084 9160
rect 5868 9120 5874 9132
rect 13078 9120 13084 9132
rect 13136 9160 13142 9172
rect 13262 9160 13268 9172
rect 13136 9132 13268 9160
rect 13136 9120 13142 9132
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 17681 9163 17739 9169
rect 17681 9160 17693 9163
rect 15160 9132 17693 9160
rect 15160 9120 15166 9132
rect 17681 9129 17693 9132
rect 17727 9129 17739 9163
rect 17681 9123 17739 9129
rect 17773 9163 17831 9169
rect 17773 9129 17785 9163
rect 17819 9160 17831 9163
rect 18046 9160 18052 9172
rect 17819 9132 18052 9160
rect 17819 9129 17831 9132
rect 17773 9123 17831 9129
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 15746 9092 15752 9104
rect 4212 9064 15752 9092
rect 4212 9052 4218 9064
rect 15746 9052 15752 9064
rect 15804 9052 15810 9104
rect 17957 9095 18015 9101
rect 17957 9092 17969 9095
rect 16316 9064 17969 9092
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 3510 9024 3516 9036
rect 3200 8996 3516 9024
rect 3200 8984 3206 8996
rect 3510 8984 3516 8996
rect 3568 9024 3574 9036
rect 4982 9024 4988 9036
rect 3568 8996 4988 9024
rect 3568 8984 3574 8996
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 6696 8996 9260 9024
rect 6696 8984 6702 8996
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1670 8956 1676 8968
rect 1544 8928 1676 8956
rect 1544 8916 1550 8928
rect 1670 8916 1676 8928
rect 1728 8956 1734 8968
rect 1949 8959 2007 8965
rect 1949 8956 1961 8959
rect 1728 8928 1961 8956
rect 1728 8916 1734 8928
rect 1949 8925 1961 8928
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8956 2191 8959
rect 2179 8928 2774 8956
rect 2179 8925 2191 8928
rect 2133 8919 2191 8925
rect 2746 8888 2774 8928
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 8570 8956 8576 8968
rect 2924 8928 8576 8956
rect 2924 8916 2930 8928
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 9137 8959 9195 8965
rect 9137 8925 9149 8959
rect 9183 8956 9195 8959
rect 9232 8956 9260 8996
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 12342 9024 12348 9036
rect 11756 8996 12348 9024
rect 11756 8984 11762 8996
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 14182 8984 14188 9036
rect 14240 9024 14246 9036
rect 15378 9024 15384 9036
rect 14240 8996 15384 9024
rect 14240 8984 14246 8996
rect 15378 8984 15384 8996
rect 15436 9024 15442 9036
rect 16316 9024 16344 9064
rect 17957 9061 17969 9064
rect 18003 9061 18015 9095
rect 17957 9055 18015 9061
rect 15436 8996 16344 9024
rect 15436 8984 15442 8996
rect 17494 8984 17500 9036
rect 17552 9024 17558 9036
rect 17865 9027 17923 9033
rect 17865 9024 17877 9027
rect 17552 8996 17877 9024
rect 17552 8984 17558 8996
rect 17865 8993 17877 8996
rect 17911 8993 17923 9027
rect 18874 9024 18880 9036
rect 17865 8987 17923 8993
rect 18156 8996 18880 9024
rect 9183 8928 9260 8956
rect 9183 8925 9195 8928
rect 9137 8919 9195 8925
rect 14734 8916 14740 8968
rect 14792 8916 14798 8968
rect 15013 8959 15071 8965
rect 15013 8925 15025 8959
rect 15059 8925 15071 8959
rect 15013 8919 15071 8925
rect 3142 8888 3148 8900
rect 2746 8860 3148 8888
rect 3142 8848 3148 8860
rect 3200 8888 3206 8900
rect 7282 8888 7288 8900
rect 3200 8860 7288 8888
rect 3200 8848 3206 8860
rect 7282 8848 7288 8860
rect 7340 8848 7346 8900
rect 8386 8848 8392 8900
rect 8444 8888 8450 8900
rect 15028 8888 15056 8919
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 17589 8959 17647 8965
rect 17589 8956 17601 8959
rect 15252 8928 17601 8956
rect 15252 8916 15258 8928
rect 17589 8925 17601 8928
rect 17635 8925 17647 8959
rect 17589 8919 17647 8925
rect 17954 8916 17960 8968
rect 18012 8916 18018 8968
rect 18156 8965 18184 8996
rect 18874 8984 18880 8996
rect 18932 8984 18938 9036
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 8444 8860 15056 8888
rect 8444 8848 8450 8860
rect 17494 8848 17500 8900
rect 17552 8888 17558 8900
rect 18248 8888 18276 8919
rect 17552 8860 18276 8888
rect 17552 8848 17558 8860
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 7064 8792 9045 8820
rect 7064 8780 7070 8792
rect 9033 8789 9045 8792
rect 9079 8789 9091 8823
rect 9033 8783 9091 8789
rect 14369 8823 14427 8829
rect 14369 8789 14381 8823
rect 14415 8820 14427 8823
rect 14642 8820 14648 8832
rect 14415 8792 14648 8820
rect 14415 8789 14427 8792
rect 14369 8783 14427 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 15010 8780 15016 8832
rect 15068 8820 15074 8832
rect 17586 8820 17592 8832
rect 15068 8792 17592 8820
rect 15068 8780 15074 8792
rect 17586 8780 17592 8792
rect 17644 8780 17650 8832
rect 18414 8780 18420 8832
rect 18472 8780 18478 8832
rect 1104 8730 18860 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 17610 8730
rect 17662 8678 17674 8730
rect 17726 8678 17738 8730
rect 17790 8678 17802 8730
rect 17854 8678 17866 8730
rect 17918 8678 18860 8730
rect 1104 8656 18860 8678
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 7101 8619 7159 8625
rect 7101 8616 7113 8619
rect 5776 8588 7113 8616
rect 5776 8576 5782 8588
rect 7101 8585 7113 8588
rect 7147 8585 7159 8619
rect 7101 8579 7159 8585
rect 7374 8576 7380 8628
rect 7432 8616 7438 8628
rect 7926 8616 7932 8628
rect 7432 8588 7932 8616
rect 7432 8576 7438 8588
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 8536 8588 9996 8616
rect 8536 8576 8542 8588
rect 4798 8508 4804 8560
rect 4856 8508 4862 8560
rect 6638 8508 6644 8560
rect 6696 8508 6702 8560
rect 9582 8548 9588 8560
rect 6932 8520 9588 8548
rect 3602 8440 3608 8492
rect 3660 8440 3666 8492
rect 3694 8440 3700 8492
rect 3752 8440 3758 8492
rect 3878 8440 3884 8492
rect 3936 8440 3942 8492
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8480 4031 8483
rect 4062 8480 4068 8492
rect 4019 8452 4068 8480
rect 4019 8449 4031 8452
rect 3973 8443 4031 8449
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4816 8480 4844 8508
rect 5166 8480 5172 8492
rect 4571 8452 5172 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 6086 8440 6092 8492
rect 6144 8480 6150 8492
rect 6546 8480 6552 8492
rect 6144 8452 6552 8480
rect 6144 8440 6150 8452
rect 6546 8440 6552 8452
rect 6604 8440 6610 8492
rect 6932 8489 6960 8520
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 9968 8548 9996 8588
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 11330 8616 11336 8628
rect 11204 8588 11336 8616
rect 11204 8576 11210 8588
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 12434 8576 12440 8628
rect 12492 8576 12498 8628
rect 14185 8619 14243 8625
rect 14185 8585 14197 8619
rect 14231 8616 14243 8619
rect 14366 8616 14372 8628
rect 14231 8588 14372 8616
rect 14231 8585 14243 8588
rect 14185 8579 14243 8585
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 14553 8619 14611 8625
rect 14553 8585 14565 8619
rect 14599 8616 14611 8619
rect 18046 8616 18052 8628
rect 14599 8588 18052 8616
rect 14599 8585 14611 8588
rect 14553 8579 14611 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 16393 8551 16451 8557
rect 16393 8548 16405 8551
rect 9968 8520 16405 8548
rect 16393 8517 16405 8520
rect 16439 8517 16451 8551
rect 16393 8511 16451 8517
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 1394 8372 1400 8424
rect 1452 8372 1458 8424
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 3050 8412 3056 8424
rect 1719 8384 3056 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4798 8412 4804 8424
rect 4479 8384 4804 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4798 8372 4804 8384
rect 4856 8412 4862 8424
rect 4982 8412 4988 8424
rect 4856 8384 4988 8412
rect 4856 8372 4862 8384
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 6748 8412 6776 8443
rect 7006 8440 7012 8492
rect 7064 8440 7070 8492
rect 7561 8483 7619 8489
rect 7116 8452 7420 8480
rect 7116 8412 7144 8452
rect 6696 8384 7144 8412
rect 7193 8415 7251 8421
rect 6696 8372 6702 8384
rect 7193 8381 7205 8415
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 3421 8347 3479 8353
rect 3421 8313 3433 8347
rect 3467 8344 3479 8347
rect 7208 8344 7236 8375
rect 7282 8372 7288 8424
rect 7340 8372 7346 8424
rect 7392 8412 7420 8452
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 7650 8480 7656 8492
rect 7607 8452 7656 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 10100 8452 10149 8480
rect 10100 8440 10106 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11514 8480 11520 8492
rect 10928 8452 11520 8480
rect 10928 8440 10934 8452
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 12360 8412 12388 8443
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 14369 8483 14427 8489
rect 14369 8449 14381 8483
rect 14415 8480 14427 8483
rect 14826 8480 14832 8492
rect 14415 8452 14832 8480
rect 14415 8449 14427 8452
rect 14369 8443 14427 8449
rect 13722 8412 13728 8424
rect 7392 8384 13728 8412
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 14108 8412 14136 8443
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 15654 8440 15660 8492
rect 15712 8480 15718 8492
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 15712 8452 16129 8480
rect 15712 8440 15718 8452
rect 16117 8449 16129 8452
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 16209 8483 16267 8489
rect 16209 8449 16221 8483
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 14458 8412 14464 8424
rect 14108 8384 14464 8412
rect 14458 8372 14464 8384
rect 14516 8412 14522 8424
rect 14734 8412 14740 8424
rect 14516 8384 14740 8412
rect 14516 8372 14522 8384
rect 14734 8372 14740 8384
rect 14792 8372 14798 8424
rect 7558 8344 7564 8356
rect 3467 8316 7236 8344
rect 7300 8316 7564 8344
rect 3467 8313 3479 8316
rect 3421 8307 3479 8313
rect 4430 8236 4436 8288
rect 4488 8236 4494 8288
rect 6365 8279 6423 8285
rect 6365 8245 6377 8279
rect 6411 8276 6423 8279
rect 6454 8276 6460 8288
rect 6411 8248 6460 8276
rect 6411 8245 6423 8248
rect 6365 8239 6423 8245
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 7300 8276 7328 8316
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 8938 8344 8944 8356
rect 7668 8316 8944 8344
rect 7248 8248 7328 8276
rect 7248 8236 7254 8248
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 7668 8276 7696 8316
rect 8938 8304 8944 8316
rect 8996 8304 9002 8356
rect 9674 8304 9680 8356
rect 9732 8304 9738 8356
rect 10502 8304 10508 8356
rect 10560 8344 10566 8356
rect 16224 8344 16252 8443
rect 10560 8316 16252 8344
rect 10560 8304 10566 8316
rect 7524 8248 7696 8276
rect 7524 8236 7530 8248
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 9861 8279 9919 8285
rect 9861 8276 9873 8279
rect 9824 8248 9873 8276
rect 9824 8236 9830 8248
rect 9861 8245 9873 8248
rect 9907 8276 9919 8279
rect 12526 8276 12532 8288
rect 9907 8248 12532 8276
rect 9907 8245 9919 8248
rect 9861 8239 9919 8245
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 16117 8279 16175 8285
rect 16117 8276 16129 8279
rect 14516 8248 16129 8276
rect 14516 8236 14522 8248
rect 16117 8245 16129 8248
rect 16163 8245 16175 8279
rect 16117 8239 16175 8245
rect 1104 8186 18860 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 11950 8186
rect 12002 8134 12014 8186
rect 12066 8134 12078 8186
rect 12130 8134 12142 8186
rect 12194 8134 12206 8186
rect 12258 8134 16950 8186
rect 17002 8134 17014 8186
rect 17066 8134 17078 8186
rect 17130 8134 17142 8186
rect 17194 8134 17206 8186
rect 17258 8134 18860 8186
rect 1104 8112 18860 8134
rect 2406 8032 2412 8084
rect 2464 8072 2470 8084
rect 2501 8075 2559 8081
rect 2501 8072 2513 8075
rect 2464 8044 2513 8072
rect 2464 8032 2470 8044
rect 2501 8041 2513 8044
rect 2547 8041 2559 8075
rect 2501 8035 2559 8041
rect 3237 8075 3295 8081
rect 3237 8041 3249 8075
rect 3283 8072 3295 8075
rect 5902 8072 5908 8084
rect 3283 8044 5908 8072
rect 3283 8041 3295 8044
rect 3237 8035 3295 8041
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7650 8072 7656 8084
rect 7248 8044 7656 8072
rect 7248 8032 7254 8044
rect 7650 8032 7656 8044
rect 7708 8072 7714 8084
rect 11514 8072 11520 8084
rect 7708 8044 11520 8072
rect 7708 8032 7714 8044
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 17865 8075 17923 8081
rect 17865 8072 17877 8075
rect 17552 8044 17877 8072
rect 17552 8032 17558 8044
rect 17865 8041 17877 8044
rect 17911 8041 17923 8075
rect 17865 8035 17923 8041
rect 3970 8004 3976 8016
rect 2056 7976 3976 8004
rect 2056 7877 2084 7976
rect 3970 7964 3976 7976
rect 4028 7964 4034 8016
rect 16298 8004 16304 8016
rect 4724 7976 16304 8004
rect 2685 7939 2743 7945
rect 2685 7905 2697 7939
rect 2731 7936 2743 7939
rect 3602 7936 3608 7948
rect 2731 7908 3608 7936
rect 2731 7905 2743 7908
rect 2685 7899 2743 7905
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 3896 7908 4660 7936
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7837 2099 7871
rect 2041 7831 2099 7837
rect 2314 7828 2320 7880
rect 2372 7828 2378 7880
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 2593 7871 2651 7877
rect 2593 7868 2605 7871
rect 2556 7840 2605 7868
rect 2556 7828 2562 7840
rect 2593 7837 2605 7840
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2958 7868 2964 7880
rect 2823 7840 2964 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 3896 7868 3924 7908
rect 3467 7840 3924 7868
rect 3973 7871 4031 7877
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4154 7868 4160 7880
rect 4019 7840 4160 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 3605 7803 3663 7809
rect 3605 7769 3617 7803
rect 3651 7800 3663 7803
rect 4246 7800 4252 7812
rect 3651 7772 4252 7800
rect 3651 7769 3663 7772
rect 3605 7763 3663 7769
rect 4246 7760 4252 7772
rect 4304 7760 4310 7812
rect 1578 7692 1584 7744
rect 1636 7732 1642 7744
rect 2133 7735 2191 7741
rect 2133 7732 2145 7735
rect 1636 7704 2145 7732
rect 1636 7692 1642 7704
rect 2133 7701 2145 7704
rect 2179 7732 2191 7735
rect 3418 7732 3424 7744
rect 2179 7704 3424 7732
rect 2179 7701 2191 7704
rect 2133 7695 2191 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 4356 7732 4384 7831
rect 4632 7800 4660 7908
rect 4724 7877 4752 7976
rect 16298 7964 16304 7976
rect 16356 7964 16362 8016
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 7098 7936 7104 7948
rect 4856 7908 7104 7936
rect 4856 7896 4862 7908
rect 7098 7896 7104 7908
rect 7156 7936 7162 7948
rect 8113 7939 8171 7945
rect 7156 7908 8064 7936
rect 7156 7896 7162 7908
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 7742 7868 7748 7880
rect 4709 7831 4767 7837
rect 4816 7840 7748 7868
rect 4816 7800 4844 7840
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 8036 7877 8064 7908
rect 8113 7905 8125 7939
rect 8159 7936 8171 7939
rect 8478 7936 8484 7948
rect 8159 7908 8484 7936
rect 8159 7905 8171 7908
rect 8113 7899 8171 7905
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 10134 7936 10140 7948
rect 8588 7908 10140 7936
rect 8588 7880 8616 7908
rect 10134 7896 10140 7908
rect 10192 7936 10198 7948
rect 14182 7936 14188 7948
rect 10192 7908 14188 7936
rect 10192 7896 10198 7908
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 8260 7840 8309 7868
rect 8260 7828 8266 7840
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7868 8447 7871
rect 8570 7868 8576 7880
rect 8435 7840 8576 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 17678 7828 17684 7880
rect 17736 7828 17742 7880
rect 4632 7772 4844 7800
rect 4893 7803 4951 7809
rect 4893 7769 4905 7803
rect 4939 7800 4951 7803
rect 9214 7800 9220 7812
rect 4939 7772 9220 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 6362 7732 6368 7744
rect 4356 7704 6368 7732
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 6638 7692 6644 7744
rect 6696 7732 6702 7744
rect 7558 7732 7564 7744
rect 6696 7704 7564 7732
rect 6696 7692 6702 7704
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 8573 7735 8631 7741
rect 8573 7732 8585 7735
rect 8352 7704 8585 7732
rect 8352 7692 8358 7704
rect 8573 7701 8585 7704
rect 8619 7701 8631 7735
rect 8573 7695 8631 7701
rect 13630 7692 13636 7744
rect 13688 7732 13694 7744
rect 14826 7732 14832 7744
rect 13688 7704 14832 7732
rect 13688 7692 13694 7704
rect 14826 7692 14832 7704
rect 14884 7732 14890 7744
rect 18966 7732 18972 7744
rect 14884 7704 18972 7732
rect 14884 7692 14890 7704
rect 18966 7692 18972 7704
rect 19024 7692 19030 7744
rect 1104 7642 18860 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 17610 7642
rect 17662 7590 17674 7642
rect 17726 7590 17738 7642
rect 17790 7590 17802 7642
rect 17854 7590 17866 7642
rect 17918 7590 18860 7642
rect 1104 7568 18860 7590
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 5258 7528 5264 7540
rect 5040 7500 5264 7528
rect 5040 7488 5046 7500
rect 5258 7488 5264 7500
rect 5316 7528 5322 7540
rect 8478 7528 8484 7540
rect 5316 7500 8484 7528
rect 5316 7488 5322 7500
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7460 1731 7463
rect 1762 7460 1768 7472
rect 1719 7432 1768 7460
rect 1719 7429 1731 7432
rect 1673 7423 1731 7429
rect 1762 7420 1768 7432
rect 1820 7420 1826 7472
rect 7098 7420 7104 7472
rect 7156 7460 7162 7472
rect 8113 7463 8171 7469
rect 8113 7460 8125 7463
rect 7156 7432 8125 7460
rect 7156 7420 7162 7432
rect 8113 7429 8125 7432
rect 8159 7429 8171 7463
rect 8113 7423 8171 7429
rect 842 7352 848 7404
rect 900 7392 906 7404
rect 1489 7395 1547 7401
rect 1489 7392 1501 7395
rect 900 7364 1501 7392
rect 900 7352 906 7364
rect 1489 7361 1501 7364
rect 1535 7361 1547 7395
rect 1489 7355 1547 7361
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7892 7364 7941 7392
rect 7892 7352 7898 7364
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 8220 7392 8248 7500
rect 8478 7488 8484 7500
rect 8536 7528 8542 7540
rect 13341 7531 13399 7537
rect 8536 7500 12434 7528
rect 8536 7488 8542 7500
rect 12406 7472 12434 7500
rect 13341 7497 13353 7531
rect 13387 7528 13399 7531
rect 13906 7528 13912 7540
rect 13387 7500 13912 7528
rect 13387 7497 13399 7500
rect 13341 7491 13399 7497
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 14369 7531 14427 7537
rect 14369 7497 14381 7531
rect 14415 7528 14427 7531
rect 16850 7528 16856 7540
rect 14415 7500 16856 7528
rect 14415 7497 14427 7500
rect 14369 7491 14427 7497
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 11422 7460 11428 7472
rect 11204 7432 11428 7460
rect 11204 7420 11210 7432
rect 11422 7420 11428 7432
rect 11480 7420 11486 7472
rect 12406 7432 12440 7472
rect 12434 7420 12440 7432
rect 12492 7420 12498 7472
rect 13541 7463 13599 7469
rect 13541 7429 13553 7463
rect 13587 7460 13599 7463
rect 13630 7460 13636 7472
rect 13587 7432 13636 7460
rect 13587 7429 13599 7432
rect 13541 7423 13599 7429
rect 13630 7420 13636 7432
rect 13688 7420 13694 7472
rect 13740 7432 16252 7460
rect 8067 7364 8248 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7392 8447 7395
rect 13740 7392 13768 7432
rect 8435 7364 13768 7392
rect 8435 7361 8447 7364
rect 8389 7355 8447 7361
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 14090 7352 14096 7404
rect 14148 7352 14154 7404
rect 14182 7352 14188 7404
rect 14240 7352 14246 7404
rect 16224 7392 16252 7432
rect 16850 7392 16856 7404
rect 16224 7364 16856 7392
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 13832 7324 13860 7352
rect 11204 7296 13860 7324
rect 13909 7327 13967 7333
rect 11204 7284 11210 7296
rect 13909 7293 13921 7327
rect 13955 7324 13967 7327
rect 13998 7324 14004 7336
rect 13955 7296 14004 7324
rect 13955 7293 13967 7296
rect 13909 7287 13967 7293
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 16298 7284 16304 7336
rect 16356 7284 16362 7336
rect 6178 7216 6184 7268
rect 6236 7256 6242 7268
rect 15933 7259 15991 7265
rect 15933 7256 15945 7259
rect 6236 7228 15945 7256
rect 6236 7216 6242 7228
rect 15933 7225 15945 7228
rect 15979 7225 15991 7259
rect 15933 7219 15991 7225
rect 1670 7148 1676 7200
rect 1728 7188 1734 7200
rect 2498 7188 2504 7200
rect 1728 7160 2504 7188
rect 1728 7148 1734 7160
rect 2498 7148 2504 7160
rect 2556 7188 2562 7200
rect 7190 7188 7196 7200
rect 2556 7160 7196 7188
rect 2556 7148 2562 7160
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 7745 7191 7803 7197
rect 7745 7188 7757 7191
rect 7524 7160 7757 7188
rect 7524 7148 7530 7160
rect 7745 7157 7757 7160
rect 7791 7157 7803 7191
rect 7745 7151 7803 7157
rect 11330 7148 11336 7200
rect 11388 7188 11394 7200
rect 13173 7191 13231 7197
rect 13173 7188 13185 7191
rect 11388 7160 13185 7188
rect 11388 7148 11394 7160
rect 13173 7157 13185 7160
rect 13219 7157 13231 7191
rect 13173 7151 13231 7157
rect 13357 7191 13415 7197
rect 13357 7157 13369 7191
rect 13403 7188 13415 7191
rect 14458 7188 14464 7200
rect 13403 7160 14464 7188
rect 13403 7157 13415 7160
rect 13357 7151 13415 7157
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 15841 7191 15899 7197
rect 15841 7188 15853 7191
rect 15252 7160 15853 7188
rect 15252 7148 15258 7160
rect 15841 7157 15853 7160
rect 15887 7157 15899 7191
rect 15841 7151 15899 7157
rect 1104 7098 18860 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 11950 7098
rect 12002 7046 12014 7098
rect 12066 7046 12078 7098
rect 12130 7046 12142 7098
rect 12194 7046 12206 7098
rect 12258 7046 16950 7098
rect 17002 7046 17014 7098
rect 17066 7046 17078 7098
rect 17130 7046 17142 7098
rect 17194 7046 17206 7098
rect 17258 7046 18860 7098
rect 1104 7024 18860 7046
rect 6546 6944 6552 6996
rect 6604 6984 6610 6996
rect 6914 6984 6920 6996
rect 6604 6956 6920 6984
rect 6604 6944 6610 6956
rect 6914 6944 6920 6956
rect 6972 6984 6978 6996
rect 7834 6984 7840 6996
rect 6972 6956 7840 6984
rect 6972 6944 6978 6956
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 9306 6944 9312 6996
rect 9364 6984 9370 6996
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 9364 6956 9413 6984
rect 9364 6944 9370 6956
rect 9401 6953 9413 6956
rect 9447 6953 9459 6987
rect 10870 6984 10876 6996
rect 9401 6947 9459 6953
rect 9508 6956 10876 6984
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 7006 6916 7012 6928
rect 4212 6888 7012 6916
rect 4212 6876 4218 6888
rect 7006 6876 7012 6888
rect 7064 6916 7070 6928
rect 9508 6916 9536 6956
rect 10870 6944 10876 6956
rect 10928 6984 10934 6996
rect 16298 6984 16304 6996
rect 10928 6956 16304 6984
rect 10928 6944 10934 6956
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 7064 6888 9536 6916
rect 12268 6888 12756 6916
rect 7064 6876 7070 6888
rect 2406 6808 2412 6860
rect 2464 6848 2470 6860
rect 2593 6851 2651 6857
rect 2593 6848 2605 6851
rect 2464 6820 2605 6848
rect 2464 6808 2470 6820
rect 2593 6817 2605 6820
rect 2639 6817 2651 6851
rect 2593 6811 2651 6817
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6848 5135 6851
rect 8386 6848 8392 6860
rect 5123 6820 8392 6848
rect 5123 6817 5135 6820
rect 5077 6811 5135 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 10134 6808 10140 6860
rect 10192 6848 10198 6860
rect 12268 6848 12296 6888
rect 10192 6820 12296 6848
rect 10192 6808 10198 6820
rect 12342 6808 12348 6860
rect 12400 6848 12406 6860
rect 12400 6820 12664 6848
rect 12400 6808 12406 6820
rect 1762 6740 1768 6792
rect 1820 6780 1826 6792
rect 2777 6783 2835 6789
rect 1820 6752 2728 6780
rect 1820 6740 1826 6752
rect 2700 6712 2728 6752
rect 2777 6749 2789 6783
rect 2823 6780 2835 6783
rect 3050 6780 3056 6792
rect 2823 6752 3056 6780
rect 2823 6749 2835 6752
rect 2777 6743 2835 6749
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4982 6780 4988 6792
rect 4212 6752 4988 6780
rect 4212 6740 4218 6752
rect 4982 6740 4988 6752
rect 5040 6740 5046 6792
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6780 5227 6783
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 5215 6752 9689 6780
rect 5215 6749 5227 6752
rect 5169 6743 5227 6749
rect 9677 6749 9689 6752
rect 9723 6780 9735 6783
rect 9766 6780 9772 6792
rect 9723 6752 9772 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 9950 6740 9956 6792
rect 10008 6740 10014 6792
rect 10042 6740 10048 6792
rect 10100 6740 10106 6792
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 12437 6783 12495 6789
rect 12437 6780 12449 6783
rect 11112 6752 12449 6780
rect 11112 6740 11118 6752
rect 12437 6749 12449 6752
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 12526 6740 12532 6792
rect 12584 6740 12590 6792
rect 12636 6789 12664 6820
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6749 12679 6783
rect 12728 6780 12756 6888
rect 16022 6876 16028 6928
rect 16080 6876 16086 6928
rect 16114 6876 16120 6928
rect 16172 6916 16178 6928
rect 16172 6888 16252 6916
rect 16172 6876 16178 6888
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 16040 6848 16068 6876
rect 16224 6857 16252 6888
rect 16209 6851 16267 6857
rect 14056 6820 15792 6848
rect 16040 6820 16160 6848
rect 14056 6808 14062 6820
rect 15764 6789 15792 6820
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 12728 6752 15301 6780
rect 12621 6743 12679 6749
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 16025 6783 16083 6789
rect 16025 6749 16037 6783
rect 16071 6749 16083 6783
rect 16132 6780 16160 6820
rect 16209 6817 16221 6851
rect 16255 6817 16267 6851
rect 16209 6811 16267 6817
rect 16132 6752 16252 6780
rect 16025 6743 16083 6749
rect 2958 6712 2964 6724
rect 2700 6684 2964 6712
rect 2958 6672 2964 6684
rect 3016 6672 3022 6724
rect 3145 6715 3203 6721
rect 3145 6681 3157 6715
rect 3191 6712 3203 6715
rect 6822 6712 6828 6724
rect 3191 6684 6828 6712
rect 3191 6681 3203 6684
rect 3145 6675 3203 6681
rect 6822 6672 6828 6684
rect 6880 6672 6886 6724
rect 8938 6672 8944 6724
rect 8996 6712 9002 6724
rect 9585 6715 9643 6721
rect 9585 6712 9597 6715
rect 8996 6684 9597 6712
rect 8996 6672 9002 6684
rect 9585 6681 9597 6684
rect 9631 6681 9643 6715
rect 9585 6675 9643 6681
rect 9861 6715 9919 6721
rect 9861 6681 9873 6715
rect 9907 6681 9919 6715
rect 10060 6712 10088 6740
rect 11146 6712 11152 6724
rect 10060 6684 11152 6712
rect 9861 6675 9919 6681
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3326 6644 3332 6656
rect 2915 6616 3332 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 5166 6604 5172 6656
rect 5224 6644 5230 6656
rect 9217 6647 9275 6653
rect 9217 6644 9229 6647
rect 5224 6616 9229 6644
rect 5224 6604 5230 6616
rect 9217 6613 9229 6616
rect 9263 6613 9275 6647
rect 9217 6607 9275 6613
rect 9385 6647 9443 6653
rect 9385 6613 9397 6647
rect 9431 6644 9443 6647
rect 9766 6644 9772 6656
rect 9431 6616 9772 6644
rect 9431 6613 9443 6616
rect 9385 6607 9443 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 9876 6644 9904 6675
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 11514 6672 11520 6724
rect 11572 6712 11578 6724
rect 12342 6712 12348 6724
rect 11572 6684 12348 6712
rect 11572 6672 11578 6684
rect 12342 6672 12348 6684
rect 12400 6672 12406 6724
rect 15654 6672 15660 6724
rect 15712 6712 15718 6724
rect 16040 6712 16068 6743
rect 16224 6724 16252 6752
rect 16758 6740 16764 6792
rect 16816 6740 16822 6792
rect 18233 6783 18291 6789
rect 18233 6749 18245 6783
rect 18279 6780 18291 6783
rect 18782 6780 18788 6792
rect 18279 6752 18788 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 15712 6684 16068 6712
rect 15712 6672 15718 6684
rect 16206 6672 16212 6724
rect 16264 6672 16270 6724
rect 9950 6644 9956 6656
rect 9876 6616 9956 6644
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10229 6647 10287 6653
rect 10229 6613 10241 6647
rect 10275 6644 10287 6647
rect 13998 6644 14004 6656
rect 10275 6616 14004 6644
rect 10275 6613 10287 6616
rect 10229 6607 10287 6613
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 18414 6604 18420 6656
rect 18472 6604 18478 6656
rect 1104 6554 18860 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 17610 6554
rect 17662 6502 17674 6554
rect 17726 6502 17738 6554
rect 17790 6502 17802 6554
rect 17854 6502 17866 6554
rect 17918 6502 18860 6554
rect 1104 6480 18860 6502
rect 2038 6400 2044 6452
rect 2096 6400 2102 6452
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 6632 6443 6690 6449
rect 6632 6440 6644 6443
rect 5868 6412 6644 6440
rect 5868 6400 5874 6412
rect 6632 6409 6644 6412
rect 6678 6440 6690 6443
rect 9674 6440 9680 6452
rect 6678 6412 9680 6440
rect 6678 6409 6690 6412
rect 6632 6403 6690 6409
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 10413 6443 10471 6449
rect 9824 6412 10272 6440
rect 9824 6400 9830 6412
rect 1394 6332 1400 6384
rect 1452 6332 1458 6384
rect 1613 6375 1671 6381
rect 1613 6341 1625 6375
rect 1659 6372 1671 6375
rect 2314 6372 2320 6384
rect 1659 6344 2320 6372
rect 1659 6341 1671 6344
rect 1613 6335 1671 6341
rect 2314 6332 2320 6344
rect 2372 6332 2378 6384
rect 2958 6332 2964 6384
rect 3016 6372 3022 6384
rect 10134 6372 10140 6384
rect 3016 6344 10140 6372
rect 3016 6332 3022 6344
rect 10134 6332 10140 6344
rect 10192 6332 10198 6384
rect 10244 6372 10272 6412
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 10594 6440 10600 6452
rect 10459 6412 10600 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 18138 6400 18144 6452
rect 18196 6440 18202 6452
rect 18233 6443 18291 6449
rect 18233 6440 18245 6443
rect 18196 6412 18245 6440
rect 18196 6400 18202 6412
rect 18233 6409 18245 6412
rect 18279 6409 18291 6443
rect 18233 6403 18291 6409
rect 10686 6372 10692 6384
rect 10244 6344 10692 6372
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 13722 6332 13728 6384
rect 13780 6332 13786 6384
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 992 6276 1869 6304
rect 992 6264 998 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 7006 6264 7012 6316
rect 7064 6264 7070 6316
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 9490 6304 9496 6316
rect 8904 6276 9496 6304
rect 8904 6264 8910 6276
rect 9490 6264 9496 6276
rect 9548 6304 9554 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9548 6276 9965 6304
rect 9548 6264 9554 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 14274 6304 14280 6316
rect 9953 6267 10011 6273
rect 10612 6276 14280 6304
rect 1394 6196 1400 6248
rect 1452 6236 1458 6248
rect 10042 6236 10048 6248
rect 1452 6208 10048 6236
rect 1452 6196 1458 6208
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 1762 6128 1768 6180
rect 1820 6128 1826 6180
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 9950 6168 9956 6180
rect 4764 6140 9956 6168
rect 4764 6128 4770 6140
rect 9950 6128 9956 6140
rect 10008 6128 10014 6180
rect 1578 6060 1584 6112
rect 1636 6060 1642 6112
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 6236 6072 6653 6100
rect 6236 6060 6242 6072
rect 6641 6069 6653 6072
rect 6687 6069 6699 6103
rect 6641 6063 6699 6069
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10612 6100 10640 6276
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 16209 6307 16267 6313
rect 16209 6273 16221 6307
rect 16255 6304 16267 6307
rect 16298 6304 16304 6316
rect 16255 6276 16304 6304
rect 16255 6273 16267 6276
rect 16209 6267 16267 6273
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 16482 6264 16488 6316
rect 16540 6304 16546 6316
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 16540 6276 18521 6304
rect 16540 6264 16546 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 12342 6236 12348 6248
rect 11848 6208 12348 6236
rect 11848 6196 11854 6208
rect 12342 6196 12348 6208
rect 12400 6236 12406 6248
rect 13265 6239 13323 6245
rect 12400 6208 13216 6236
rect 12400 6196 12406 6208
rect 10284 6072 10640 6100
rect 10284 6060 10290 6072
rect 10686 6060 10692 6112
rect 10744 6100 10750 6112
rect 12434 6100 12440 6112
rect 10744 6072 12440 6100
rect 10744 6060 10750 6072
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 13188 6100 13216 6208
rect 13265 6205 13277 6239
rect 13311 6236 13323 6239
rect 13814 6236 13820 6248
rect 13311 6208 13820 6236
rect 13311 6205 13323 6208
rect 13265 6199 13323 6205
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 16114 6196 16120 6248
rect 16172 6196 16178 6248
rect 18230 6196 18236 6248
rect 18288 6196 18294 6248
rect 13354 6128 13360 6180
rect 13412 6128 13418 6180
rect 15838 6128 15844 6180
rect 15896 6128 15902 6180
rect 16206 6128 16212 6180
rect 16264 6168 16270 6180
rect 16482 6168 16488 6180
rect 16264 6140 16488 6168
rect 16264 6128 16270 6140
rect 16482 6128 16488 6140
rect 16540 6128 16546 6180
rect 16758 6128 16764 6180
rect 16816 6168 16822 6180
rect 18417 6171 18475 6177
rect 18417 6168 18429 6171
rect 16816 6140 18429 6168
rect 16816 6128 16822 6140
rect 18417 6137 18429 6140
rect 18463 6137 18475 6171
rect 18417 6131 18475 6137
rect 18322 6100 18328 6112
rect 13188 6072 18328 6100
rect 18322 6060 18328 6072
rect 18380 6060 18386 6112
rect 1104 6010 18860 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 11950 6010
rect 12002 5958 12014 6010
rect 12066 5958 12078 6010
rect 12130 5958 12142 6010
rect 12194 5958 12206 6010
rect 12258 5958 16950 6010
rect 17002 5958 17014 6010
rect 17066 5958 17078 6010
rect 17130 5958 17142 6010
rect 17194 5958 17206 6010
rect 17258 5958 18860 6010
rect 1104 5936 18860 5958
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 3234 5896 3240 5908
rect 2372 5868 3240 5896
rect 2372 5856 2378 5868
rect 3234 5856 3240 5868
rect 3292 5896 3298 5908
rect 4062 5896 4068 5908
rect 3292 5868 4068 5896
rect 3292 5856 3298 5868
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5865 4307 5899
rect 4249 5859 4307 5865
rect 4264 5828 4292 5859
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4396 5868 4445 5896
rect 4396 5856 4402 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 6638 5856 6644 5908
rect 6696 5896 6702 5908
rect 6696 5868 11928 5896
rect 6696 5856 6702 5868
rect 4706 5828 4712 5840
rect 4264 5800 4712 5828
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 11900 5828 11928 5868
rect 13170 5856 13176 5908
rect 13228 5896 13234 5908
rect 14737 5899 14795 5905
rect 13228 5868 14688 5896
rect 13228 5856 13234 5868
rect 13814 5828 13820 5840
rect 8168 5800 11652 5828
rect 11900 5800 13820 5828
rect 8168 5788 8174 5800
rect 11422 5720 11428 5772
rect 11480 5760 11486 5772
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 11480 5732 11529 5760
rect 11480 5720 11486 5732
rect 11517 5729 11529 5732
rect 11563 5729 11575 5763
rect 11624 5760 11652 5800
rect 13814 5788 13820 5800
rect 13872 5788 13878 5840
rect 14093 5763 14151 5769
rect 14093 5760 14105 5763
rect 11624 5732 14105 5760
rect 11517 5723 11575 5729
rect 4522 5692 4528 5704
rect 4080 5664 4528 5692
rect 4080 5633 4108 5664
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 12176 5701 12204 5732
rect 14093 5729 14105 5732
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 11885 5695 11943 5701
rect 11885 5692 11897 5695
rect 10928 5664 11897 5692
rect 10928 5652 10934 5664
rect 11885 5661 11897 5664
rect 11931 5661 11943 5695
rect 11885 5655 11943 5661
rect 12161 5695 12219 5701
rect 12161 5661 12173 5695
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 4065 5627 4123 5633
rect 4065 5593 4077 5627
rect 4111 5593 4123 5627
rect 4065 5587 4123 5593
rect 4281 5627 4339 5633
rect 4281 5593 4293 5627
rect 4327 5624 4339 5627
rect 9306 5624 9312 5636
rect 4327 5596 9312 5624
rect 4327 5593 4339 5596
rect 4281 5587 4339 5593
rect 9306 5584 9312 5596
rect 9364 5584 9370 5636
rect 11900 5556 11928 5655
rect 12342 5652 12348 5704
rect 12400 5692 12406 5704
rect 12897 5695 12955 5701
rect 12897 5692 12909 5695
rect 12400 5664 12909 5692
rect 12400 5652 12406 5664
rect 12897 5661 12909 5664
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 13449 5695 13507 5701
rect 13449 5661 13461 5695
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 13464 5624 13492 5655
rect 13538 5652 13544 5704
rect 13596 5692 13602 5704
rect 14185 5695 14243 5701
rect 14185 5692 14197 5695
rect 13596 5664 14197 5692
rect 13596 5652 13602 5664
rect 14185 5661 14197 5664
rect 14231 5661 14243 5695
rect 14185 5655 14243 5661
rect 14274 5652 14280 5704
rect 14332 5692 14338 5704
rect 14660 5701 14688 5868
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 14826 5896 14832 5908
rect 14783 5868 14832 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 14826 5856 14832 5868
rect 14884 5896 14890 5908
rect 15010 5896 15016 5908
rect 14884 5868 15016 5896
rect 14884 5856 14890 5868
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 16574 5856 16580 5908
rect 16632 5896 16638 5908
rect 16761 5899 16819 5905
rect 16761 5896 16773 5899
rect 16632 5868 16773 5896
rect 16632 5856 16638 5868
rect 16761 5865 16773 5868
rect 16807 5865 16819 5899
rect 16761 5859 16819 5865
rect 15930 5720 15936 5772
rect 15988 5760 15994 5772
rect 15988 5732 16436 5760
rect 15988 5720 15994 5732
rect 14369 5695 14427 5701
rect 14369 5692 14381 5695
rect 14332 5664 14381 5692
rect 14332 5652 14338 5664
rect 14369 5661 14381 5664
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 14826 5652 14832 5704
rect 14884 5652 14890 5704
rect 15378 5652 15384 5704
rect 15436 5692 15442 5704
rect 16408 5701 16436 5732
rect 16482 5720 16488 5772
rect 16540 5760 16546 5772
rect 16540 5732 16896 5760
rect 16540 5720 16546 5732
rect 16868 5701 16896 5732
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 15436 5664 16129 5692
rect 15436 5652 15442 5664
rect 16117 5661 16129 5664
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5661 16451 5695
rect 16393 5655 16451 5661
rect 16853 5695 16911 5701
rect 16853 5661 16865 5695
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 16482 5624 16488 5636
rect 13096 5596 13308 5624
rect 13464 5596 16488 5624
rect 13096 5556 13124 5596
rect 11900 5528 13124 5556
rect 13170 5516 13176 5568
rect 13228 5516 13234 5568
rect 13280 5556 13308 5596
rect 16482 5584 16488 5596
rect 16540 5584 16546 5636
rect 16577 5627 16635 5633
rect 16577 5593 16589 5627
rect 16623 5624 16635 5627
rect 18230 5624 18236 5636
rect 16623 5596 18236 5624
rect 16623 5593 16635 5596
rect 16577 5587 16635 5593
rect 18230 5584 18236 5596
rect 18288 5584 18294 5636
rect 13538 5556 13544 5568
rect 13280 5528 13544 5556
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 14550 5516 14556 5568
rect 14608 5516 14614 5568
rect 16206 5516 16212 5568
rect 16264 5516 16270 5568
rect 1104 5466 18860 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 17610 5466
rect 17662 5414 17674 5466
rect 17726 5414 17738 5466
rect 17790 5414 17802 5466
rect 17854 5414 17866 5466
rect 17918 5414 18860 5466
rect 1104 5392 18860 5414
rect 1486 5312 1492 5364
rect 1544 5352 1550 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1544 5324 1593 5352
rect 1544 5312 1550 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 4154 5352 4160 5364
rect 2547 5324 4160 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 5261 5355 5319 5361
rect 5261 5321 5273 5355
rect 5307 5352 5319 5355
rect 7374 5352 7380 5364
rect 5307 5324 7380 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 8018 5312 8024 5364
rect 8076 5312 8082 5364
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 15381 5355 15439 5361
rect 11112 5324 14688 5352
rect 11112 5312 11118 5324
rect 7837 5287 7895 5293
rect 7837 5284 7849 5287
rect 7392 5256 7849 5284
rect 7392 5228 7420 5256
rect 7837 5253 7849 5256
rect 7883 5284 7895 5287
rect 10870 5284 10876 5296
rect 7883 5256 10876 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 11977 5287 12035 5293
rect 11977 5253 11989 5287
rect 12023 5284 12035 5287
rect 12023 5256 12848 5284
rect 12023 5253 12035 5256
rect 11977 5247 12035 5253
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 6822 5216 6828 5228
rect 2271 5188 6828 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 7374 5176 7380 5228
rect 7432 5176 7438 5228
rect 7742 5176 7748 5228
rect 7800 5176 7806 5228
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5216 8171 5219
rect 8159 5188 8248 5216
rect 8159 5185 8171 5188
rect 8113 5179 8171 5185
rect 4801 5151 4859 5157
rect 4801 5117 4813 5151
rect 4847 5148 4859 5151
rect 7929 5151 7987 5157
rect 4847 5120 7880 5148
rect 4847 5117 4859 5120
rect 4801 5111 4859 5117
rect 5166 5040 5172 5092
rect 5224 5040 5230 5092
rect 6914 5040 6920 5092
rect 6972 5080 6978 5092
rect 7742 5080 7748 5092
rect 6972 5052 7748 5080
rect 6972 5040 6978 5052
rect 7742 5040 7748 5052
rect 7800 5040 7806 5092
rect 7852 5080 7880 5120
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 8018 5148 8024 5160
rect 7975 5120 8024 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 8220 5148 8248 5188
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 11992 5216 12020 5247
rect 8352 5188 12020 5216
rect 8352 5176 8358 5188
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12820 5225 12848 5256
rect 12986 5244 12992 5296
rect 13044 5244 13050 5296
rect 14550 5284 14556 5296
rect 13096 5256 14556 5284
rect 12621 5219 12679 5225
rect 12621 5216 12633 5219
rect 12308 5188 12633 5216
rect 12308 5176 12314 5188
rect 12621 5185 12633 5188
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 12805 5219 12863 5225
rect 12805 5185 12817 5219
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 13096 5148 13124 5256
rect 14550 5244 14556 5256
rect 14608 5244 14614 5296
rect 14660 5284 14688 5324
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 16206 5352 16212 5364
rect 15427 5324 16212 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 16390 5284 16396 5296
rect 14660 5256 16396 5284
rect 16390 5244 16396 5256
rect 16448 5244 16454 5296
rect 13262 5176 13268 5228
rect 13320 5216 13326 5228
rect 13357 5219 13415 5225
rect 13357 5216 13369 5219
rect 13320 5188 13369 5216
rect 13320 5176 13326 5188
rect 13357 5185 13369 5188
rect 13403 5185 13415 5219
rect 13357 5179 13415 5185
rect 13446 5176 13452 5228
rect 13504 5176 13510 5228
rect 13722 5176 13728 5228
rect 13780 5176 13786 5228
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5216 15255 5219
rect 15286 5216 15292 5228
rect 15243 5188 15292 5216
rect 15243 5185 15255 5188
rect 15197 5179 15255 5185
rect 15286 5176 15292 5188
rect 15344 5176 15350 5228
rect 15378 5176 15384 5228
rect 15436 5176 15442 5228
rect 8220 5120 13124 5148
rect 13170 5108 13176 5160
rect 13228 5108 13234 5160
rect 11054 5080 11060 5092
rect 7852 5052 11060 5080
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 11698 5040 11704 5092
rect 11756 5080 11762 5092
rect 11756 5052 12434 5080
rect 11756 5040 11762 5052
rect 3050 4972 3056 5024
rect 3108 5012 3114 5024
rect 8294 5012 8300 5024
rect 3108 4984 8300 5012
rect 3108 4972 3114 4984
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 9306 5012 9312 5024
rect 9088 4984 9312 5012
rect 9088 4972 9094 4984
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 11146 4972 11152 5024
rect 11204 5012 11210 5024
rect 11422 5012 11428 5024
rect 11204 4984 11428 5012
rect 11204 4972 11210 4984
rect 11422 4972 11428 4984
rect 11480 5012 11486 5024
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 11480 4984 12081 5012
rect 11480 4972 11486 4984
rect 12069 4981 12081 4984
rect 12115 4981 12127 5015
rect 12406 5012 12434 5052
rect 13633 5015 13691 5021
rect 13633 5012 13645 5015
rect 12406 4984 13645 5012
rect 12069 4975 12127 4981
rect 13633 4981 13645 4984
rect 13679 5012 13691 5015
rect 16758 5012 16764 5024
rect 13679 4984 16764 5012
rect 13679 4981 13691 4984
rect 13633 4975 13691 4981
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 1104 4922 18860 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 11950 4922
rect 12002 4870 12014 4922
rect 12066 4870 12078 4922
rect 12130 4870 12142 4922
rect 12194 4870 12206 4922
rect 12258 4870 16950 4922
rect 17002 4870 17014 4922
rect 17066 4870 17078 4922
rect 17130 4870 17142 4922
rect 17194 4870 17206 4922
rect 17258 4870 18860 4922
rect 1104 4848 18860 4870
rect 13722 4808 13728 4820
rect 2746 4780 13728 4808
rect 1486 4700 1492 4752
rect 1544 4740 1550 4752
rect 2746 4740 2774 4780
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14090 4768 14096 4820
rect 14148 4768 14154 4820
rect 14277 4811 14335 4817
rect 14277 4808 14289 4811
rect 14200 4780 14289 4808
rect 1544 4712 2774 4740
rect 1544 4700 1550 4712
rect 4062 4700 4068 4752
rect 4120 4740 4126 4752
rect 10045 4743 10103 4749
rect 10045 4740 10057 4743
rect 4120 4712 10057 4740
rect 4120 4700 4126 4712
rect 10045 4709 10057 4712
rect 10091 4709 10103 4743
rect 10045 4703 10103 4709
rect 12066 4700 12072 4752
rect 12124 4700 12130 4752
rect 12434 4700 12440 4752
rect 12492 4700 12498 4752
rect 13078 4700 13084 4752
rect 13136 4740 13142 4752
rect 14200 4740 14228 4780
rect 14277 4777 14289 4780
rect 14323 4777 14335 4811
rect 16298 4808 16304 4820
rect 14277 4771 14335 4777
rect 16040 4780 16304 4808
rect 13136 4712 14228 4740
rect 13136 4700 13142 4712
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 8938 4672 8944 4684
rect 6880 4644 8944 4672
rect 6880 4632 6886 4644
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 9214 4632 9220 4684
rect 9272 4632 9278 4684
rect 9306 4632 9312 4684
rect 9364 4632 9370 4684
rect 9401 4675 9459 4681
rect 9401 4641 9413 4675
rect 9447 4672 9459 4675
rect 10226 4672 10232 4684
rect 9447 4644 10232 4672
rect 9447 4641 9459 4644
rect 9401 4635 9459 4641
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 12526 4632 12532 4684
rect 12584 4632 12590 4684
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 16040 4672 16068 4780
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 16666 4768 16672 4820
rect 16724 4768 16730 4820
rect 16761 4811 16819 4817
rect 16761 4777 16773 4811
rect 16807 4808 16819 4811
rect 16850 4808 16856 4820
rect 16807 4780 16856 4808
rect 16807 4777 16819 4780
rect 16761 4771 16819 4777
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 18506 4740 18512 4752
rect 13872 4644 16068 4672
rect 16132 4712 18512 4740
rect 13872 4632 13878 4644
rect 8846 4564 8852 4616
rect 8904 4604 8910 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 8904 4576 9137 4604
rect 8904 4564 8910 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 9030 4536 9036 4548
rect 7800 4508 9036 4536
rect 7800 4496 7806 4508
rect 9030 4496 9036 4508
rect 9088 4496 9094 4548
rect 10888 4536 10916 4567
rect 11054 4564 11060 4616
rect 11112 4564 11118 4616
rect 11606 4564 11612 4616
rect 11664 4604 11670 4616
rect 12253 4607 12311 4613
rect 12253 4604 12265 4607
rect 11664 4576 12265 4604
rect 11664 4564 11670 4576
rect 12253 4573 12265 4576
rect 12299 4573 12311 4607
rect 12253 4567 12311 4573
rect 14458 4564 14464 4616
rect 14516 4604 14522 4616
rect 14645 4607 14703 4613
rect 14645 4604 14657 4607
rect 14516 4576 14657 4604
rect 14516 4564 14522 4576
rect 14645 4573 14657 4576
rect 14691 4573 14703 4607
rect 14645 4567 14703 4573
rect 15654 4564 15660 4616
rect 15712 4604 15718 4616
rect 16132 4613 16160 4712
rect 18506 4700 18512 4712
rect 18564 4700 18570 4752
rect 16025 4607 16083 4613
rect 16025 4604 16037 4607
rect 15712 4576 16037 4604
rect 15712 4564 15718 4576
rect 16025 4573 16037 4576
rect 16071 4573 16083 4607
rect 16025 4567 16083 4573
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4573 16175 4607
rect 16485 4607 16543 4613
rect 16485 4604 16497 4607
rect 16117 4567 16175 4573
rect 16224 4576 16497 4604
rect 11146 4536 11152 4548
rect 10888 4508 11152 4536
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 11992 4508 12204 4536
rect 8938 4428 8944 4480
rect 8996 4428 9002 4480
rect 9306 4428 9312 4480
rect 9364 4468 9370 4480
rect 11992 4468 12020 4508
rect 9364 4440 12020 4468
rect 12176 4468 12204 4508
rect 12342 4496 12348 4548
rect 12400 4536 12406 4548
rect 16224 4536 16252 4576
rect 16485 4573 16497 4576
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 16758 4564 16764 4616
rect 16816 4564 16822 4616
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 12400 4508 16252 4536
rect 12400 4496 12406 4508
rect 16298 4496 16304 4548
rect 16356 4496 16362 4548
rect 16390 4496 16396 4548
rect 16448 4496 16454 4548
rect 13814 4468 13820 4480
rect 12176 4440 13820 4468
rect 9364 4428 9370 4440
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 13998 4428 14004 4480
rect 14056 4468 14062 4480
rect 14277 4471 14335 4477
rect 14277 4468 14289 4471
rect 14056 4440 14289 4468
rect 14056 4428 14062 4440
rect 14277 4437 14289 4440
rect 14323 4437 14335 4471
rect 14277 4431 14335 4437
rect 14918 4428 14924 4480
rect 14976 4468 14982 4480
rect 16960 4468 16988 4567
rect 14976 4440 16988 4468
rect 14976 4428 14982 4440
rect 1104 4378 18860 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 17610 4378
rect 17662 4326 17674 4378
rect 17726 4326 17738 4378
rect 17790 4326 17802 4378
rect 17854 4326 17866 4378
rect 17918 4326 18860 4378
rect 1104 4304 18860 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 9306 4264 9312 4276
rect 2464 4236 9312 4264
rect 2464 4224 2470 4236
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 9858 4224 9864 4276
rect 9916 4264 9922 4276
rect 10045 4267 10103 4273
rect 10045 4264 10057 4267
rect 9916 4236 10057 4264
rect 9916 4224 9922 4236
rect 10045 4233 10057 4236
rect 10091 4233 10103 4267
rect 10045 4227 10103 4233
rect 10134 4224 10140 4276
rect 10192 4224 10198 4276
rect 3142 4156 3148 4208
rect 3200 4156 3206 4208
rect 9950 4156 9956 4208
rect 10008 4196 10014 4208
rect 10229 4199 10287 4205
rect 10229 4196 10241 4199
rect 10008 4168 10241 4196
rect 10008 4156 10014 4168
rect 10229 4165 10241 4168
rect 10275 4165 10287 4199
rect 10229 4159 10287 4165
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 14521 4199 14579 4205
rect 14521 4196 14533 4199
rect 11112 4168 14533 4196
rect 11112 4156 11118 4168
rect 14521 4165 14533 4168
rect 14567 4165 14579 4199
rect 14521 4159 14579 4165
rect 14734 4156 14740 4208
rect 14792 4156 14798 4208
rect 15102 4156 15108 4208
rect 15160 4196 15166 4208
rect 16390 4196 16396 4208
rect 15160 4168 16396 4196
rect 15160 4156 15166 4168
rect 16390 4156 16396 4168
rect 16448 4156 16454 4208
rect 17494 4156 17500 4208
rect 17552 4196 17558 4208
rect 17954 4196 17960 4208
rect 17552 4168 17960 4196
rect 17552 4156 17558 4168
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 900 4100 1409 4128
rect 900 4088 906 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 5644 4060 5672 4091
rect 5810 4088 5816 4140
rect 5868 4088 5874 4140
rect 8754 4088 8760 4140
rect 8812 4128 8818 4140
rect 10134 4128 10140 4140
rect 8812 4100 10140 4128
rect 8812 4088 8818 4100
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 15194 4128 15200 4140
rect 12360 4100 15200 4128
rect 12360 4060 12388 4100
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 15286 4088 15292 4140
rect 15344 4128 15350 4140
rect 17313 4131 17371 4137
rect 17313 4128 17325 4131
rect 15344 4100 17325 4128
rect 15344 4088 15350 4100
rect 17313 4097 17325 4100
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 18230 4088 18236 4140
rect 18288 4088 18294 4140
rect 5644 4032 12388 4060
rect 17681 4063 17739 4069
rect 17681 4029 17693 4063
rect 17727 4060 17739 4063
rect 18322 4060 18328 4072
rect 17727 4032 18328 4060
rect 17727 4029 17739 4032
rect 17681 4023 17739 4029
rect 18322 4020 18328 4032
rect 18380 4020 18386 4072
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 1854 3992 1860 4004
rect 1627 3964 1860 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 1854 3952 1860 3964
rect 1912 3952 1918 4004
rect 5810 3952 5816 4004
rect 5868 3952 5874 4004
rect 9861 3995 9919 4001
rect 9861 3961 9873 3995
rect 9907 3992 9919 3995
rect 10318 3992 10324 4004
rect 9907 3964 10324 3992
rect 9907 3961 9919 3964
rect 9861 3955 9919 3961
rect 10318 3952 10324 3964
rect 10376 3952 10382 4004
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 12400 3964 14596 3992
rect 12400 3952 12406 3964
rect 3053 3927 3111 3933
rect 3053 3893 3065 3927
rect 3099 3924 3111 3927
rect 3234 3924 3240 3936
rect 3099 3896 3240 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 10413 3927 10471 3933
rect 10413 3924 10425 3927
rect 9456 3896 10425 3924
rect 9456 3884 9462 3896
rect 10413 3893 10425 3896
rect 10459 3893 10471 3927
rect 10413 3887 10471 3893
rect 14366 3884 14372 3936
rect 14424 3884 14430 3936
rect 14568 3933 14596 3964
rect 14553 3927 14611 3933
rect 14553 3893 14565 3927
rect 14599 3924 14611 3927
rect 16206 3924 16212 3936
rect 14599 3896 16212 3924
rect 14599 3893 14611 3896
rect 14553 3887 14611 3893
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 18414 3884 18420 3936
rect 18472 3884 18478 3936
rect 1104 3834 18860 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 11950 3834
rect 12002 3782 12014 3834
rect 12066 3782 12078 3834
rect 12130 3782 12142 3834
rect 12194 3782 12206 3834
rect 12258 3782 16950 3834
rect 17002 3782 17014 3834
rect 17066 3782 17078 3834
rect 17130 3782 17142 3834
rect 17194 3782 17206 3834
rect 17258 3782 18860 3834
rect 1104 3760 18860 3782
rect 3878 3680 3884 3732
rect 3936 3680 3942 3732
rect 4341 3723 4399 3729
rect 4341 3689 4353 3723
rect 4387 3720 4399 3723
rect 7282 3720 7288 3732
rect 4387 3692 7288 3720
rect 4387 3689 4399 3692
rect 4341 3683 4399 3689
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 15102 3720 15108 3732
rect 9416 3692 15108 3720
rect 5074 3612 5080 3664
rect 5132 3652 5138 3664
rect 9125 3655 9183 3661
rect 9125 3652 9137 3655
rect 5132 3624 9137 3652
rect 5132 3612 5138 3624
rect 9125 3621 9137 3624
rect 9171 3621 9183 3655
rect 9125 3615 9183 3621
rect 1854 3544 1860 3596
rect 1912 3584 1918 3596
rect 9416 3584 9444 3692
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 15289 3723 15347 3729
rect 15289 3689 15301 3723
rect 15335 3720 15347 3723
rect 17310 3720 17316 3732
rect 15335 3692 17316 3720
rect 15335 3689 15347 3692
rect 15289 3683 15347 3689
rect 17310 3680 17316 3692
rect 17368 3680 17374 3732
rect 13446 3652 13452 3664
rect 1912 3556 9444 3584
rect 1912 3544 1918 3556
rect 3602 3476 3608 3528
rect 3660 3516 3666 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3660 3488 3801 3516
rect 3660 3476 3666 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4080 3448 4108 3479
rect 9306 3476 9312 3528
rect 9364 3476 9370 3528
rect 9416 3525 9444 3556
rect 9508 3624 13452 3652
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 4246 3448 4252 3460
rect 4080 3420 4252 3448
rect 4246 3408 4252 3420
rect 4304 3448 4310 3460
rect 9125 3451 9183 3457
rect 9125 3448 9137 3451
rect 4304 3420 9137 3448
rect 4304 3408 4310 3420
rect 9125 3417 9137 3420
rect 9171 3448 9183 3451
rect 9508 3448 9536 3624
rect 13446 3612 13452 3624
rect 13504 3612 13510 3664
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 14458 3584 14464 3596
rect 11204 3556 14464 3584
rect 11204 3544 11210 3556
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3584 14703 3587
rect 15470 3584 15476 3596
rect 14691 3556 15476 3584
rect 14691 3553 14703 3556
rect 14645 3547 14703 3553
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 11330 3516 11336 3528
rect 9640 3488 11336 3516
rect 9640 3476 9646 3488
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 13078 3516 13084 3528
rect 12216 3488 13084 3516
rect 12216 3476 12222 3488
rect 13078 3476 13084 3488
rect 13136 3516 13142 3528
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 13136 3488 15025 3516
rect 13136 3476 13142 3488
rect 15013 3485 15025 3488
rect 15059 3485 15071 3519
rect 15013 3479 15071 3485
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3485 15163 3519
rect 15105 3479 15163 3485
rect 9171 3420 9536 3448
rect 9171 3417 9183 3420
rect 9125 3411 9183 3417
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 15120 3448 15148 3479
rect 11296 3420 15148 3448
rect 11296 3408 11302 3420
rect 10962 3340 10968 3392
rect 11020 3380 11026 3392
rect 12526 3380 12532 3392
rect 11020 3352 12532 3380
rect 11020 3340 11026 3352
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 1104 3290 18860 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 17610 3290
rect 17662 3238 17674 3290
rect 17726 3238 17738 3290
rect 17790 3238 17802 3290
rect 17854 3238 17866 3290
rect 17918 3238 18860 3290
rect 1104 3216 18860 3238
rect 9582 3176 9588 3188
rect 2746 3148 9588 3176
rect 1670 3068 1676 3120
rect 1728 3068 1734 3120
rect 842 3000 848 3052
rect 900 3040 906 3052
rect 1489 3043 1547 3049
rect 1489 3040 1501 3043
rect 900 3012 1501 3040
rect 900 3000 906 3012
rect 1489 3009 1501 3012
rect 1535 3009 1547 3043
rect 1489 3003 1547 3009
rect 1854 3000 1860 3052
rect 1912 3000 1918 3052
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 2746 3040 2774 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 11020 3148 12296 3176
rect 11020 3136 11026 3148
rect 3970 3108 3976 3120
rect 3804 3080 3976 3108
rect 3804 3049 3832 3080
rect 3970 3068 3976 3080
rect 4028 3068 4034 3120
rect 4065 3111 4123 3117
rect 4065 3077 4077 3111
rect 4111 3108 4123 3111
rect 4246 3108 4252 3120
rect 4111 3080 4252 3108
rect 4111 3077 4123 3080
rect 4065 3071 4123 3077
rect 4246 3068 4252 3080
rect 4304 3068 4310 3120
rect 6454 3068 6460 3120
rect 6512 3108 6518 3120
rect 12268 3117 12296 3148
rect 12253 3111 12311 3117
rect 6512 3080 12020 3108
rect 6512 3068 6518 3080
rect 2363 3012 2774 3040
rect 3789 3043 3847 3049
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 3789 3009 3801 3043
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 4798 3040 4804 3052
rect 3927 3012 4804 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 2148 2972 2176 3003
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8904 3012 8953 3040
rect 8904 3000 8910 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3009 9183 3043
rect 9125 3003 9183 3009
rect 9140 2972 9168 3003
rect 9214 3000 9220 3052
rect 9272 3000 9278 3052
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 10686 3040 10692 3052
rect 10560 3012 10692 3040
rect 10560 3000 10566 3012
rect 10686 3000 10692 3012
rect 10744 3040 10750 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10744 3012 10977 3040
rect 10744 3000 10750 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11146 3000 11152 3052
rect 11204 3000 11210 3052
rect 11422 3040 11428 3052
rect 11256 3012 11428 3040
rect 11256 2972 11284 3012
rect 11422 3000 11428 3012
rect 11480 3000 11486 3052
rect 11992 3049 12020 3080
rect 12253 3077 12265 3111
rect 12299 3077 12311 3111
rect 12253 3071 12311 3077
rect 12342 3068 12348 3120
rect 12400 3068 12406 3120
rect 13906 3068 13912 3120
rect 13964 3108 13970 3120
rect 14277 3111 14335 3117
rect 14277 3108 14289 3111
rect 13964 3080 14289 3108
rect 13964 3068 13970 3080
rect 14277 3077 14289 3080
rect 14323 3077 14335 3111
rect 14277 3071 14335 3077
rect 14461 3111 14519 3117
rect 14461 3077 14473 3111
rect 14507 3108 14519 3111
rect 15010 3108 15016 3120
rect 14507 3080 15016 3108
rect 14507 3077 14519 3080
rect 14461 3071 14519 3077
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 12158 3049 12164 3052
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12125 3043 12164 3049
rect 12125 3009 12137 3043
rect 12125 3003 12164 3009
rect 12158 3000 12164 3003
rect 12216 3000 12222 3052
rect 12526 3049 12532 3052
rect 12483 3043 12532 3049
rect 12483 3009 12495 3043
rect 12529 3009 12532 3043
rect 12483 3003 12532 3009
rect 12526 3000 12532 3003
rect 12584 3000 12590 3052
rect 14550 3000 14556 3052
rect 14608 3000 14614 3052
rect 2148 2944 7604 2972
rect 9140 2944 11284 2972
rect 11333 2975 11391 2981
rect 2041 2907 2099 2913
rect 2041 2873 2053 2907
rect 2087 2904 2099 2907
rect 7374 2904 7380 2916
rect 2087 2876 7380 2904
rect 2087 2873 2099 2876
rect 2041 2867 2099 2873
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 7576 2904 7604 2944
rect 11333 2941 11345 2975
rect 11379 2972 11391 2975
rect 14642 2972 14648 2984
rect 11379 2944 14648 2972
rect 11379 2941 11391 2944
rect 11333 2935 11391 2941
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 14277 2907 14335 2913
rect 14277 2904 14289 2907
rect 7576 2876 14289 2904
rect 14277 2873 14289 2876
rect 14323 2873 14335 2907
rect 14277 2867 14335 2873
rect 2314 2796 2320 2848
rect 2372 2796 2378 2848
rect 4065 2839 4123 2845
rect 4065 2805 4077 2839
rect 4111 2836 4123 2839
rect 8202 2836 8208 2848
rect 4111 2808 8208 2836
rect 4111 2805 4123 2808
rect 4065 2799 4123 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 12621 2839 12679 2845
rect 12621 2805 12633 2839
rect 12667 2836 12679 2839
rect 18690 2836 18696 2848
rect 12667 2808 18696 2836
rect 12667 2805 12679 2808
rect 12621 2799 12679 2805
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 1104 2746 18860 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 11950 2746
rect 12002 2694 12014 2746
rect 12066 2694 12078 2746
rect 12130 2694 12142 2746
rect 12194 2694 12206 2746
rect 12258 2694 16950 2746
rect 17002 2694 17014 2746
rect 17066 2694 17078 2746
rect 17130 2694 17142 2746
rect 17194 2694 17206 2746
rect 17258 2694 18860 2746
rect 1104 2672 18860 2694
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4614 2632 4620 2644
rect 4203 2604 4620 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2632 9091 2635
rect 11054 2632 11060 2644
rect 9079 2604 11060 2632
rect 9079 2601 9091 2604
rect 9033 2595 9091 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 15562 2592 15568 2644
rect 15620 2632 15626 2644
rect 17865 2635 17923 2641
rect 17865 2632 17877 2635
rect 15620 2604 17877 2632
rect 15620 2592 15626 2604
rect 17865 2601 17877 2604
rect 17911 2601 17923 2635
rect 17865 2595 17923 2601
rect 1302 2524 1308 2576
rect 1360 2564 1366 2576
rect 1857 2567 1915 2573
rect 1857 2564 1869 2567
rect 1360 2536 1869 2564
rect 1360 2524 1366 2536
rect 1857 2533 1869 2536
rect 1903 2533 1915 2567
rect 1857 2527 1915 2533
rect 10413 2567 10471 2573
rect 10413 2533 10425 2567
rect 10459 2564 10471 2567
rect 10778 2564 10784 2576
rect 10459 2536 10784 2564
rect 10459 2533 10471 2536
rect 10413 2527 10471 2533
rect 10778 2524 10784 2536
rect 10836 2564 10842 2576
rect 15286 2564 15292 2576
rect 10836 2536 15292 2564
rect 10836 2524 10842 2536
rect 15286 2524 15292 2536
rect 15344 2524 15350 2576
rect 17402 2524 17408 2576
rect 17460 2564 17466 2576
rect 17681 2567 17739 2573
rect 17681 2564 17693 2567
rect 17460 2536 17693 2564
rect 17460 2524 17466 2536
rect 17681 2533 17693 2536
rect 17727 2533 17739 2567
rect 17681 2527 17739 2533
rect 10686 2496 10692 2508
rect 1688 2468 10692 2496
rect 1688 2437 1716 2468
rect 10686 2456 10692 2468
rect 10744 2456 10750 2508
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 17494 2496 17500 2508
rect 16991 2468 17500 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 7466 2428 7472 2440
rect 2363 2400 7472 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 1780 2360 1808 2391
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 8938 2388 8944 2440
rect 8996 2388 9002 2440
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 15746 2388 15752 2440
rect 15804 2388 15810 2440
rect 16574 2388 16580 2440
rect 16632 2428 16638 2440
rect 16761 2431 16819 2437
rect 16761 2428 16773 2431
rect 16632 2400 16773 2428
rect 16632 2388 16638 2400
rect 16761 2397 16773 2400
rect 16807 2397 16819 2431
rect 16761 2391 16819 2397
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18598 2428 18604 2440
rect 18279 2400 18604 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 1268 2332 1808 2360
rect 1268 2320 1274 2332
rect 3326 2320 3332 2372
rect 3384 2360 3390 2372
rect 3881 2363 3939 2369
rect 3881 2360 3893 2363
rect 3384 2332 3893 2360
rect 3384 2320 3390 2332
rect 3881 2329 3893 2332
rect 3927 2329 3939 2363
rect 3881 2323 3939 2329
rect 9950 2320 9956 2372
rect 10008 2360 10014 2372
rect 10137 2363 10195 2369
rect 10137 2360 10149 2363
rect 10008 2332 10149 2360
rect 10008 2320 10014 2332
rect 10137 2329 10149 2332
rect 10183 2329 10195 2363
rect 10137 2323 10195 2329
rect 13722 2320 13728 2372
rect 13780 2360 13786 2372
rect 15933 2363 15991 2369
rect 15933 2360 15945 2363
rect 13780 2332 15945 2360
rect 13780 2320 13786 2332
rect 15933 2329 15945 2332
rect 15979 2329 15991 2363
rect 15933 2323 15991 2329
rect 16114 2320 16120 2372
rect 16172 2320 16178 2372
rect 16206 2320 16212 2372
rect 16264 2360 16270 2372
rect 17833 2363 17891 2369
rect 17833 2360 17845 2363
rect 16264 2332 17845 2360
rect 16264 2320 16270 2332
rect 17833 2329 17845 2332
rect 17879 2329 17891 2363
rect 17833 2323 17891 2329
rect 18046 2320 18052 2372
rect 18104 2320 18110 2372
rect 18414 2252 18420 2304
rect 18472 2252 18478 2304
rect 1104 2202 18860 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 17610 2202
rect 17662 2150 17674 2202
rect 17726 2150 17738 2202
rect 17790 2150 17802 2202
rect 17854 2150 17866 2202
rect 17918 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 5448 17620 5500 17672
rect 18144 17620 18196 17672
rect 13268 17552 13320 17604
rect 16580 17552 16632 17604
rect 9312 17484 9364 17536
rect 18236 17484 18288 17536
rect 2610 17382 2662 17434
rect 2674 17382 2726 17434
rect 2738 17382 2790 17434
rect 2802 17382 2854 17434
rect 2866 17382 2918 17434
rect 7610 17382 7662 17434
rect 7674 17382 7726 17434
rect 7738 17382 7790 17434
rect 7802 17382 7854 17434
rect 7866 17382 7918 17434
rect 12610 17382 12662 17434
rect 12674 17382 12726 17434
rect 12738 17382 12790 17434
rect 12802 17382 12854 17434
rect 12866 17382 12918 17434
rect 17610 17382 17662 17434
rect 17674 17382 17726 17434
rect 17738 17382 17790 17434
rect 17802 17382 17854 17434
rect 17866 17382 17918 17434
rect 1860 17255 1912 17264
rect 1860 17221 1869 17255
rect 1869 17221 1903 17255
rect 1903 17221 1912 17255
rect 1860 17212 1912 17221
rect 13268 17280 13320 17332
rect 17960 17280 18012 17332
rect 848 17144 900 17196
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 5080 17144 5132 17196
rect 10508 17212 10560 17264
rect 13636 17212 13688 17264
rect 13728 17212 13780 17264
rect 8852 17144 8904 17196
rect 2320 17008 2372 17060
rect 1400 16940 1452 16992
rect 10048 17076 10100 17128
rect 14464 17076 14516 17128
rect 15200 17119 15252 17128
rect 15200 17085 15209 17119
rect 15209 17085 15243 17119
rect 15243 17085 15252 17119
rect 15200 17076 15252 17085
rect 16396 17144 16448 17196
rect 18236 17187 18288 17196
rect 18236 17153 18245 17187
rect 18245 17153 18279 17187
rect 18279 17153 18288 17187
rect 18236 17144 18288 17153
rect 4160 17008 4212 17060
rect 10232 17008 10284 17060
rect 11796 17008 11848 17060
rect 15660 17008 15712 17060
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5540 16940 5592 16992
rect 9772 16940 9824 16992
rect 10784 16940 10836 16992
rect 14648 16940 14700 16992
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 6950 16838 7002 16890
rect 7014 16838 7066 16890
rect 7078 16838 7130 16890
rect 7142 16838 7194 16890
rect 7206 16838 7258 16890
rect 11950 16838 12002 16890
rect 12014 16838 12066 16890
rect 12078 16838 12130 16890
rect 12142 16838 12194 16890
rect 12206 16838 12258 16890
rect 16950 16838 17002 16890
rect 17014 16838 17066 16890
rect 17078 16838 17130 16890
rect 17142 16838 17194 16890
rect 17206 16838 17258 16890
rect 4988 16736 5040 16788
rect 5448 16736 5500 16788
rect 4160 16711 4212 16720
rect 4160 16677 4169 16711
rect 4169 16677 4203 16711
rect 4203 16677 4212 16711
rect 4160 16668 4212 16677
rect 5540 16575 5592 16584
rect 5540 16541 5549 16575
rect 5549 16541 5583 16575
rect 5583 16541 5592 16575
rect 5540 16532 5592 16541
rect 8300 16736 8352 16788
rect 9496 16736 9548 16788
rect 9864 16736 9916 16788
rect 6552 16668 6604 16720
rect 3700 16464 3752 16516
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 9680 16668 9732 16720
rect 11244 16736 11296 16788
rect 15660 16779 15712 16788
rect 15660 16745 15669 16779
rect 15669 16745 15703 16779
rect 15703 16745 15712 16779
rect 15660 16736 15712 16745
rect 6736 16575 6788 16584
rect 6736 16541 6745 16575
rect 6745 16541 6779 16575
rect 6779 16541 6788 16575
rect 6736 16532 6788 16541
rect 8392 16532 8444 16584
rect 8760 16532 8812 16584
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 9588 16532 9640 16584
rect 10048 16532 10100 16584
rect 10324 16575 10376 16584
rect 10324 16541 10333 16575
rect 10333 16541 10367 16575
rect 10367 16541 10376 16575
rect 10324 16532 10376 16541
rect 13912 16668 13964 16720
rect 10692 16600 10744 16652
rect 13636 16600 13688 16652
rect 14280 16600 14332 16652
rect 10876 16532 10928 16584
rect 7380 16464 7432 16516
rect 9956 16507 10008 16516
rect 9956 16473 9965 16507
rect 9965 16473 9999 16507
rect 9999 16473 10008 16507
rect 9956 16464 10008 16473
rect 10600 16507 10652 16516
rect 10600 16473 10609 16507
rect 10609 16473 10643 16507
rect 10643 16473 10652 16507
rect 10600 16464 10652 16473
rect 12440 16464 12492 16516
rect 14464 16575 14516 16584
rect 14464 16541 14473 16575
rect 14473 16541 14507 16575
rect 14507 16541 14516 16575
rect 14464 16532 14516 16541
rect 14648 16643 14700 16652
rect 14648 16609 14657 16643
rect 14657 16609 14691 16643
rect 14691 16609 14700 16643
rect 14648 16600 14700 16609
rect 16764 16668 16816 16720
rect 18328 16736 18380 16788
rect 18512 16668 18564 16720
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 15200 16575 15252 16584
rect 15200 16541 15209 16575
rect 15209 16541 15243 16575
rect 15243 16541 15252 16575
rect 15200 16532 15252 16541
rect 13268 16464 13320 16516
rect 14188 16507 14240 16516
rect 14188 16473 14197 16507
rect 14197 16473 14231 16507
rect 14231 16473 14240 16507
rect 14188 16464 14240 16473
rect 7288 16396 7340 16448
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 10140 16396 10192 16448
rect 10324 16396 10376 16448
rect 11152 16396 11204 16448
rect 14924 16396 14976 16448
rect 15384 16464 15436 16516
rect 16672 16532 16724 16584
rect 18788 16600 18840 16652
rect 16856 16575 16908 16584
rect 16856 16541 16865 16575
rect 16865 16541 16899 16575
rect 16899 16541 16908 16575
rect 16856 16532 16908 16541
rect 16948 16532 17000 16584
rect 17316 16464 17368 16516
rect 17408 16464 17460 16516
rect 15936 16396 15988 16448
rect 17500 16396 17552 16448
rect 17960 16439 18012 16448
rect 17960 16405 17969 16439
rect 17969 16405 18003 16439
rect 18003 16405 18012 16439
rect 17960 16396 18012 16405
rect 18420 16396 18472 16448
rect 2610 16294 2662 16346
rect 2674 16294 2726 16346
rect 2738 16294 2790 16346
rect 2802 16294 2854 16346
rect 2866 16294 2918 16346
rect 7610 16294 7662 16346
rect 7674 16294 7726 16346
rect 7738 16294 7790 16346
rect 7802 16294 7854 16346
rect 7866 16294 7918 16346
rect 12610 16294 12662 16346
rect 12674 16294 12726 16346
rect 12738 16294 12790 16346
rect 12802 16294 12854 16346
rect 12866 16294 12918 16346
rect 17610 16294 17662 16346
rect 17674 16294 17726 16346
rect 17738 16294 17790 16346
rect 17802 16294 17854 16346
rect 17866 16294 17918 16346
rect 2964 16192 3016 16244
rect 5632 16192 5684 16244
rect 9496 16192 9548 16244
rect 11520 16192 11572 16244
rect 13176 16192 13228 16244
rect 15476 16192 15528 16244
rect 1032 16124 1084 16176
rect 1584 16056 1636 16108
rect 2504 16056 2556 16108
rect 4068 16124 4120 16176
rect 9404 16124 9456 16176
rect 9864 16124 9916 16176
rect 3056 16099 3108 16108
rect 3056 16065 3065 16099
rect 3065 16065 3099 16099
rect 3099 16065 3108 16099
rect 3056 16056 3108 16065
rect 3148 16056 3200 16108
rect 9956 16056 10008 16108
rect 10048 16056 10100 16108
rect 11980 16124 12032 16176
rect 18880 16124 18932 16176
rect 12992 16056 13044 16108
rect 13268 16056 13320 16108
rect 13452 16056 13504 16108
rect 14556 16056 14608 16108
rect 18144 16056 18196 16108
rect 18604 16056 18656 16108
rect 4804 15988 4856 16040
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 1492 15963 1544 15972
rect 1492 15929 1501 15963
rect 1501 15929 1535 15963
rect 1535 15929 1544 15963
rect 1492 15920 1544 15929
rect 9220 15920 9272 15972
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 10968 15988 11020 16040
rect 11336 15988 11388 16040
rect 12900 15988 12952 16040
rect 14924 15988 14976 16040
rect 11428 15920 11480 15972
rect 15476 15920 15528 15972
rect 9864 15895 9916 15904
rect 9864 15861 9873 15895
rect 9873 15861 9907 15895
rect 9907 15861 9916 15895
rect 9864 15852 9916 15861
rect 11060 15852 11112 15904
rect 11796 15852 11848 15904
rect 14648 15852 14700 15904
rect 15844 15852 15896 15904
rect 17960 15852 18012 15904
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 6950 15750 7002 15802
rect 7014 15750 7066 15802
rect 7078 15750 7130 15802
rect 7142 15750 7194 15802
rect 7206 15750 7258 15802
rect 11950 15750 12002 15802
rect 12014 15750 12066 15802
rect 12078 15750 12130 15802
rect 12142 15750 12194 15802
rect 12206 15750 12258 15802
rect 16950 15750 17002 15802
rect 17014 15750 17066 15802
rect 17078 15750 17130 15802
rect 17142 15750 17194 15802
rect 17206 15750 17258 15802
rect 10968 15648 11020 15700
rect 11428 15648 11480 15700
rect 14096 15648 14148 15700
rect 5724 15580 5776 15632
rect 2412 15512 2464 15564
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 8484 15512 8536 15564
rect 10692 15512 10744 15564
rect 10968 15555 11020 15564
rect 10968 15521 10977 15555
rect 10977 15521 11011 15555
rect 11011 15521 11020 15555
rect 10968 15512 11020 15521
rect 13544 15555 13596 15564
rect 13544 15521 13553 15555
rect 13553 15521 13587 15555
rect 13587 15521 13596 15555
rect 13544 15512 13596 15521
rect 13728 15512 13780 15564
rect 2964 15376 3016 15428
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 10416 15444 10468 15496
rect 13176 15444 13228 15496
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 14924 15444 14976 15496
rect 15476 15487 15528 15496
rect 15476 15453 15485 15487
rect 15485 15453 15519 15487
rect 15519 15453 15528 15487
rect 15476 15444 15528 15453
rect 16580 15444 16632 15496
rect 17132 15487 17184 15496
rect 17132 15453 17141 15487
rect 17141 15453 17175 15487
rect 17175 15453 17184 15487
rect 17132 15444 17184 15453
rect 18052 15444 18104 15496
rect 18144 15444 18196 15496
rect 5816 15308 5868 15360
rect 6368 15308 6420 15360
rect 12900 15376 12952 15428
rect 13268 15376 13320 15428
rect 8116 15308 8168 15360
rect 9036 15308 9088 15360
rect 15384 15376 15436 15428
rect 16856 15419 16908 15428
rect 16856 15385 16865 15419
rect 16865 15385 16899 15419
rect 16899 15385 16908 15419
rect 16856 15376 16908 15385
rect 17960 15308 18012 15360
rect 18696 15376 18748 15428
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 7610 15206 7662 15258
rect 7674 15206 7726 15258
rect 7738 15206 7790 15258
rect 7802 15206 7854 15258
rect 7866 15206 7918 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 17610 15206 17662 15258
rect 17674 15206 17726 15258
rect 17738 15206 17790 15258
rect 17802 15206 17854 15258
rect 17866 15206 17918 15258
rect 3884 15104 3936 15156
rect 8944 15104 8996 15156
rect 9680 15104 9732 15156
rect 848 14968 900 15020
rect 5540 15036 5592 15088
rect 3516 15011 3568 15020
rect 3516 14977 3525 15011
rect 3525 14977 3559 15011
rect 3559 14977 3568 15011
rect 3516 14968 3568 14977
rect 6644 14968 6696 15020
rect 7656 15011 7708 15020
rect 7656 14977 7665 15011
rect 7665 14977 7699 15011
rect 7699 14977 7708 15011
rect 7656 14968 7708 14977
rect 8576 15036 8628 15088
rect 9404 15036 9456 15088
rect 10692 15104 10744 15156
rect 3424 14764 3476 14816
rect 7472 14900 7524 14952
rect 8208 14968 8260 15020
rect 6736 14832 6788 14884
rect 6092 14764 6144 14816
rect 7564 14764 7616 14816
rect 8024 14832 8076 14884
rect 8668 14832 8720 14884
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 10600 14968 10652 15020
rect 12624 15036 12676 15088
rect 13728 15036 13780 15088
rect 11612 14968 11664 15020
rect 17868 15104 17920 15156
rect 18328 15104 18380 15156
rect 17132 15036 17184 15088
rect 17960 15036 18012 15088
rect 14188 14968 14240 15020
rect 14556 14968 14608 15020
rect 16120 14968 16172 15020
rect 9404 14943 9456 14952
rect 9404 14909 9413 14943
rect 9413 14909 9447 14943
rect 9447 14909 9456 14943
rect 9404 14900 9456 14909
rect 9772 14900 9824 14952
rect 9680 14832 9732 14884
rect 10140 14943 10192 14952
rect 10140 14909 10148 14943
rect 10148 14909 10182 14943
rect 10182 14909 10192 14943
rect 10140 14900 10192 14909
rect 12900 14900 12952 14952
rect 14096 14900 14148 14952
rect 14372 14900 14424 14952
rect 16764 14900 16816 14952
rect 18328 14968 18380 15020
rect 18604 14968 18656 15020
rect 17500 14900 17552 14952
rect 10508 14832 10560 14884
rect 14832 14875 14884 14884
rect 14832 14841 14841 14875
rect 14841 14841 14875 14875
rect 14875 14841 14884 14875
rect 14832 14832 14884 14841
rect 8944 14764 8996 14816
rect 9496 14807 9548 14816
rect 9496 14773 9505 14807
rect 9505 14773 9539 14807
rect 9539 14773 9548 14807
rect 9496 14764 9548 14773
rect 13544 14764 13596 14816
rect 14464 14764 14516 14816
rect 14740 14807 14792 14816
rect 14740 14773 14749 14807
rect 14749 14773 14783 14807
rect 14783 14773 14792 14807
rect 14740 14764 14792 14773
rect 16580 14764 16632 14816
rect 18880 14764 18932 14816
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 6950 14662 7002 14714
rect 7014 14662 7066 14714
rect 7078 14662 7130 14714
rect 7142 14662 7194 14714
rect 7206 14662 7258 14714
rect 11950 14662 12002 14714
rect 12014 14662 12066 14714
rect 12078 14662 12130 14714
rect 12142 14662 12194 14714
rect 12206 14662 12258 14714
rect 16950 14662 17002 14714
rect 17014 14662 17066 14714
rect 17078 14662 17130 14714
rect 17142 14662 17194 14714
rect 17206 14662 17258 14714
rect 1860 14560 1912 14612
rect 7656 14560 7708 14612
rect 9680 14560 9732 14612
rect 10140 14603 10192 14612
rect 10140 14569 10149 14603
rect 10149 14569 10183 14603
rect 10183 14569 10192 14603
rect 10140 14560 10192 14569
rect 12624 14560 12676 14612
rect 13544 14560 13596 14612
rect 14924 14560 14976 14612
rect 4160 14492 4212 14544
rect 8300 14492 8352 14544
rect 8576 14492 8628 14544
rect 12900 14492 12952 14544
rect 13084 14492 13136 14544
rect 13452 14492 13504 14544
rect 14096 14492 14148 14544
rect 7564 14424 7616 14476
rect 10232 14424 10284 14476
rect 10508 14424 10560 14476
rect 13360 14424 13412 14476
rect 15752 14424 15804 14476
rect 8116 14356 8168 14408
rect 18420 14424 18472 14476
rect 5908 14288 5960 14340
rect 8024 14220 8076 14272
rect 11704 14288 11756 14340
rect 9588 14263 9640 14272
rect 9588 14229 9597 14263
rect 9597 14229 9631 14263
rect 9631 14229 9640 14263
rect 9588 14220 9640 14229
rect 10968 14220 11020 14272
rect 14924 14220 14976 14272
rect 16764 14288 16816 14340
rect 17868 14356 17920 14408
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 17040 14263 17092 14272
rect 17040 14229 17049 14263
rect 17049 14229 17083 14263
rect 17083 14229 17092 14263
rect 17040 14220 17092 14229
rect 17408 14220 17460 14272
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 7610 14118 7662 14170
rect 7674 14118 7726 14170
rect 7738 14118 7790 14170
rect 7802 14118 7854 14170
rect 7866 14118 7918 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 17610 14118 17662 14170
rect 17674 14118 17726 14170
rect 17738 14118 17790 14170
rect 17802 14118 17854 14170
rect 17866 14118 17918 14170
rect 7564 14016 7616 14068
rect 8208 14016 8260 14068
rect 8024 13948 8076 14000
rect 8668 13948 8720 14000
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 5264 13880 5316 13932
rect 9312 14016 9364 14068
rect 9404 14016 9456 14068
rect 9588 14016 9640 14068
rect 10232 14016 10284 14068
rect 12348 13948 12400 14000
rect 12532 13948 12584 14000
rect 13360 13948 13412 14000
rect 3424 13812 3476 13864
rect 6184 13812 6236 13864
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 9128 13880 9180 13932
rect 10048 13880 10100 13932
rect 14372 13880 14424 13932
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 18420 14059 18472 14068
rect 18420 14025 18429 14059
rect 18429 14025 18463 14059
rect 18463 14025 18472 14059
rect 18420 14016 18472 14025
rect 14832 13923 14884 13932
rect 14832 13889 14841 13923
rect 14841 13889 14875 13923
rect 14875 13889 14884 13923
rect 14832 13880 14884 13889
rect 15292 13880 15344 13932
rect 8668 13812 8720 13864
rect 11428 13812 11480 13864
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 14004 13812 14056 13864
rect 14924 13812 14976 13864
rect 1676 13744 1728 13796
rect 6920 13744 6972 13796
rect 8208 13744 8260 13796
rect 8392 13744 8444 13796
rect 15108 13744 15160 13796
rect 15568 13744 15620 13796
rect 1768 13676 1820 13728
rect 6460 13676 6512 13728
rect 8116 13676 8168 13728
rect 9036 13676 9088 13728
rect 11520 13676 11572 13728
rect 12532 13676 12584 13728
rect 13544 13676 13596 13728
rect 15476 13676 15528 13728
rect 18144 13676 18196 13728
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 11950 13574 12002 13626
rect 12014 13574 12066 13626
rect 12078 13574 12130 13626
rect 12142 13574 12194 13626
rect 12206 13574 12258 13626
rect 16950 13574 17002 13626
rect 17014 13574 17066 13626
rect 17078 13574 17130 13626
rect 17142 13574 17194 13626
rect 17206 13574 17258 13626
rect 6644 13472 6696 13524
rect 7196 13472 7248 13524
rect 7932 13472 7984 13524
rect 8116 13472 8168 13524
rect 10048 13472 10100 13524
rect 5540 13404 5592 13456
rect 8944 13404 8996 13456
rect 10784 13404 10836 13456
rect 13176 13515 13228 13524
rect 13176 13481 13185 13515
rect 13185 13481 13219 13515
rect 13219 13481 13228 13515
rect 13176 13472 13228 13481
rect 13544 13472 13596 13524
rect 13820 13404 13872 13456
rect 3792 13336 3844 13388
rect 10968 13336 11020 13388
rect 11428 13336 11480 13388
rect 12256 13336 12308 13388
rect 13360 13336 13412 13388
rect 14096 13336 14148 13388
rect 2964 13268 3016 13320
rect 3332 13311 3384 13320
rect 3332 13277 3341 13311
rect 3341 13277 3375 13311
rect 3375 13277 3384 13311
rect 3332 13268 3384 13277
rect 5724 13268 5776 13320
rect 9036 13268 9088 13320
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 9404 13268 9456 13320
rect 9772 13268 9824 13320
rect 12532 13268 12584 13320
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 13728 13268 13780 13320
rect 17500 13472 17552 13524
rect 15200 13404 15252 13456
rect 15660 13336 15712 13388
rect 16212 13336 16264 13388
rect 14556 13311 14608 13320
rect 14556 13277 14565 13311
rect 14565 13277 14599 13311
rect 14599 13277 14608 13311
rect 14556 13268 14608 13277
rect 14832 13268 14884 13320
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15568 13268 15620 13277
rect 16028 13268 16080 13320
rect 3608 13200 3660 13252
rect 3976 13200 4028 13252
rect 9588 13200 9640 13252
rect 14464 13200 14516 13252
rect 4528 13132 4580 13184
rect 8392 13132 8444 13184
rect 8760 13132 8812 13184
rect 10968 13132 11020 13184
rect 14096 13132 14148 13184
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 7610 13030 7662 13082
rect 7674 13030 7726 13082
rect 7738 13030 7790 13082
rect 7802 13030 7854 13082
rect 7866 13030 7918 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 17610 13030 17662 13082
rect 17674 13030 17726 13082
rect 17738 13030 17790 13082
rect 17802 13030 17854 13082
rect 17866 13030 17918 13082
rect 1492 12928 1544 12980
rect 1860 12928 1912 12980
rect 5908 12928 5960 12980
rect 10324 12928 10376 12980
rect 10416 12928 10468 12980
rect 13084 12928 13136 12980
rect 13268 12928 13320 12980
rect 13636 12928 13688 12980
rect 14280 12928 14332 12980
rect 14556 12928 14608 12980
rect 14372 12860 14424 12912
rect 17500 12860 17552 12912
rect 848 12792 900 12844
rect 3424 12792 3476 12844
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 4436 12792 4488 12844
rect 4528 12835 4580 12844
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 5632 12792 5684 12844
rect 5724 12835 5776 12844
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 5724 12792 5776 12801
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 7472 12792 7524 12844
rect 7840 12792 7892 12844
rect 8208 12792 8260 12844
rect 8300 12835 8352 12844
rect 8300 12801 8309 12835
rect 8309 12801 8343 12835
rect 8343 12801 8352 12835
rect 8300 12792 8352 12801
rect 8852 12792 8904 12844
rect 9588 12792 9640 12844
rect 10324 12792 10376 12844
rect 5724 12656 5776 12708
rect 7288 12656 7340 12708
rect 8760 12724 8812 12776
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 10692 12792 10744 12844
rect 11796 12792 11848 12844
rect 12256 12792 12308 12844
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 14924 12792 14976 12844
rect 16764 12724 16816 12776
rect 7932 12656 7984 12708
rect 8392 12656 8444 12708
rect 11428 12656 11480 12708
rect 7380 12588 7432 12640
rect 7748 12631 7800 12640
rect 7748 12597 7757 12631
rect 7757 12597 7791 12631
rect 7791 12597 7800 12631
rect 7748 12588 7800 12597
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 8668 12588 8720 12640
rect 12992 12656 13044 12708
rect 14280 12656 14332 12708
rect 12532 12588 12584 12640
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 11950 12486 12002 12538
rect 12014 12486 12066 12538
rect 12078 12486 12130 12538
rect 12142 12486 12194 12538
rect 12206 12486 12258 12538
rect 16950 12486 17002 12538
rect 17014 12486 17066 12538
rect 17078 12486 17130 12538
rect 17142 12486 17194 12538
rect 17206 12486 17258 12538
rect 1584 12384 1636 12436
rect 1768 12316 1820 12368
rect 6736 12316 6788 12368
rect 8116 12384 8168 12436
rect 8300 12316 8352 12368
rect 2320 12180 2372 12232
rect 3332 12180 3384 12232
rect 6460 12180 6512 12232
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 7656 12180 7708 12232
rect 8024 12180 8076 12232
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 9680 12384 9732 12436
rect 10140 12384 10192 12436
rect 10416 12384 10468 12436
rect 11244 12384 11296 12436
rect 11704 12384 11756 12436
rect 11888 12384 11940 12436
rect 12992 12316 13044 12368
rect 15476 12384 15528 12436
rect 16304 12384 16356 12436
rect 16580 12384 16632 12436
rect 15200 12316 15252 12368
rect 8760 12248 8812 12300
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 11428 12248 11480 12300
rect 11888 12248 11940 12300
rect 12348 12248 12400 12300
rect 13912 12248 13964 12300
rect 14096 12248 14148 12300
rect 14372 12291 14424 12300
rect 14372 12257 14381 12291
rect 14381 12257 14415 12291
rect 14415 12257 14424 12291
rect 14372 12248 14424 12257
rect 9404 12223 9456 12232
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 4620 12112 4672 12164
rect 7196 12112 7248 12164
rect 7840 12112 7892 12164
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 11612 12180 11664 12232
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 9864 12112 9916 12164
rect 10692 12155 10744 12164
rect 10692 12121 10701 12155
rect 10701 12121 10735 12155
rect 10735 12121 10744 12155
rect 10692 12112 10744 12121
rect 12164 12223 12216 12232
rect 12164 12189 12173 12223
rect 12173 12189 12207 12223
rect 12207 12189 12216 12223
rect 12164 12180 12216 12189
rect 12624 12180 12676 12232
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 1860 12044 1912 12096
rect 6000 12044 6052 12096
rect 7564 12044 7616 12096
rect 8208 12044 8260 12096
rect 8668 12087 8720 12096
rect 8668 12053 8677 12087
rect 8677 12053 8711 12087
rect 8711 12053 8720 12087
rect 8668 12044 8720 12053
rect 9496 12044 9548 12096
rect 9680 12044 9732 12096
rect 10508 12044 10560 12096
rect 11060 12044 11112 12096
rect 11428 12044 11480 12096
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 18052 12180 18104 12232
rect 15476 12112 15528 12164
rect 13452 12044 13504 12096
rect 13912 12044 13964 12096
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 7610 11942 7662 11994
rect 7674 11942 7726 11994
rect 7738 11942 7790 11994
rect 7802 11942 7854 11994
rect 7866 11942 7918 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 17610 11942 17662 11994
rect 17674 11942 17726 11994
rect 17738 11942 17790 11994
rect 17802 11942 17854 11994
rect 17866 11942 17918 11994
rect 4252 11840 4304 11892
rect 7288 11840 7340 11892
rect 3792 11772 3844 11824
rect 6184 11772 6236 11824
rect 12716 11840 12768 11892
rect 13084 11840 13136 11892
rect 14096 11840 14148 11892
rect 15384 11840 15436 11892
rect 18696 11840 18748 11892
rect 18972 11840 19024 11892
rect 848 11704 900 11756
rect 5816 11704 5868 11756
rect 5908 11704 5960 11756
rect 6460 11704 6512 11756
rect 4068 11636 4120 11688
rect 7288 11747 7340 11756
rect 7288 11713 7297 11747
rect 7297 11713 7331 11747
rect 7331 11713 7340 11747
rect 7288 11704 7340 11713
rect 7840 11772 7892 11824
rect 9588 11772 9640 11824
rect 7564 11636 7616 11688
rect 2964 11568 3016 11620
rect 10600 11704 10652 11756
rect 7748 11636 7800 11688
rect 8484 11636 8536 11688
rect 10232 11679 10284 11688
rect 10232 11645 10241 11679
rect 10241 11645 10275 11679
rect 10275 11645 10284 11679
rect 10232 11636 10284 11645
rect 11980 11815 12032 11824
rect 11980 11781 11989 11815
rect 11989 11781 12023 11815
rect 12023 11781 12032 11815
rect 11980 11772 12032 11781
rect 11888 11704 11940 11756
rect 13176 11772 13228 11824
rect 13636 11772 13688 11824
rect 14280 11815 14332 11824
rect 14280 11781 14289 11815
rect 14289 11781 14323 11815
rect 14323 11781 14332 11815
rect 14280 11772 14332 11781
rect 14188 11704 14240 11756
rect 14556 11772 14608 11824
rect 15108 11772 15160 11824
rect 15384 11704 15436 11756
rect 18696 11704 18748 11756
rect 8208 11568 8260 11620
rect 11612 11568 11664 11620
rect 12164 11568 12216 11620
rect 15844 11636 15896 11688
rect 17316 11636 17368 11688
rect 14832 11568 14884 11620
rect 15016 11568 15068 11620
rect 18144 11636 18196 11688
rect 18604 11568 18656 11620
rect 1492 11500 1544 11552
rect 2320 11500 2372 11552
rect 3976 11543 4028 11552
rect 3976 11509 3985 11543
rect 3985 11509 4019 11543
rect 4019 11509 4028 11543
rect 3976 11500 4028 11509
rect 5816 11500 5868 11552
rect 6552 11500 6604 11552
rect 7104 11500 7156 11552
rect 7564 11500 7616 11552
rect 7656 11543 7708 11552
rect 7656 11509 7665 11543
rect 7665 11509 7699 11543
rect 7699 11509 7708 11543
rect 7656 11500 7708 11509
rect 8852 11500 8904 11552
rect 10968 11500 11020 11552
rect 11520 11500 11572 11552
rect 12072 11500 12124 11552
rect 12624 11500 12676 11552
rect 12992 11500 13044 11552
rect 13268 11500 13320 11552
rect 14372 11500 14424 11552
rect 16120 11500 16172 11552
rect 18420 11543 18472 11552
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 18420 11500 18472 11509
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 11950 11398 12002 11450
rect 12014 11398 12066 11450
rect 12078 11398 12130 11450
rect 12142 11398 12194 11450
rect 12206 11398 12258 11450
rect 16950 11398 17002 11450
rect 17014 11398 17066 11450
rect 17078 11398 17130 11450
rect 17142 11398 17194 11450
rect 17206 11398 17258 11450
rect 3332 11296 3384 11348
rect 1492 11228 1544 11280
rect 1676 11228 1728 11280
rect 3792 11228 3844 11280
rect 1676 11092 1728 11144
rect 5540 11228 5592 11280
rect 4712 11160 4764 11212
rect 5908 11339 5960 11348
rect 5908 11305 5917 11339
rect 5917 11305 5951 11339
rect 5951 11305 5960 11339
rect 5908 11296 5960 11305
rect 6460 11296 6512 11348
rect 7288 11296 7340 11348
rect 8852 11296 8904 11348
rect 9036 11296 9088 11348
rect 9220 11296 9272 11348
rect 7656 11228 7708 11280
rect 4436 11135 4488 11144
rect 4436 11101 4445 11135
rect 4445 11101 4479 11135
rect 4479 11101 4488 11135
rect 4436 11092 4488 11101
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 4344 11024 4396 11076
rect 3976 10956 4028 11008
rect 5724 11092 5776 11144
rect 7472 11160 7524 11212
rect 5356 11067 5408 11076
rect 5356 11033 5365 11067
rect 5365 11033 5399 11067
rect 5399 11033 5408 11067
rect 5356 11024 5408 11033
rect 9864 11092 9916 11144
rect 11060 11092 11112 11144
rect 11520 11092 11572 11144
rect 11796 11092 11848 11144
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 12532 11203 12584 11212
rect 12532 11169 12541 11203
rect 12541 11169 12575 11203
rect 12575 11169 12584 11203
rect 12532 11160 12584 11169
rect 14556 11228 14608 11280
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 16212 11296 16264 11348
rect 14832 11203 14884 11212
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 15568 11228 15620 11280
rect 15016 11203 15068 11212
rect 15016 11169 15025 11203
rect 15025 11169 15059 11203
rect 15059 11169 15068 11203
rect 15016 11160 15068 11169
rect 15936 11160 15988 11212
rect 14188 11092 14240 11144
rect 10876 11024 10928 11076
rect 14648 11024 14700 11076
rect 14832 11024 14884 11076
rect 6092 10956 6144 11008
rect 6460 10956 6512 11008
rect 12624 10956 12676 11008
rect 13268 10956 13320 11008
rect 14096 10956 14148 11008
rect 14464 10956 14516 11008
rect 16120 11067 16172 11076
rect 16120 11033 16129 11067
rect 16129 11033 16163 11067
rect 16163 11033 16172 11067
rect 16120 11024 16172 11033
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 17610 10854 17662 10906
rect 17674 10854 17726 10906
rect 17738 10854 17790 10906
rect 17802 10854 17854 10906
rect 17866 10854 17918 10906
rect 3976 10752 4028 10804
rect 4160 10752 4212 10804
rect 1584 10684 1636 10736
rect 3792 10727 3844 10736
rect 3792 10693 3801 10727
rect 3801 10693 3835 10727
rect 3835 10693 3844 10727
rect 3792 10684 3844 10693
rect 4528 10752 4580 10804
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 1860 10616 1912 10668
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 3516 10616 3568 10668
rect 3976 10659 4028 10668
rect 3976 10625 3985 10659
rect 3985 10625 4019 10659
rect 4019 10625 4028 10659
rect 3976 10616 4028 10625
rect 4620 10684 4672 10736
rect 4988 10795 5040 10804
rect 4988 10761 4997 10795
rect 4997 10761 5031 10795
rect 5031 10761 5040 10795
rect 4988 10752 5040 10761
rect 5356 10752 5408 10804
rect 9036 10752 9088 10804
rect 9128 10752 9180 10804
rect 15108 10752 15160 10804
rect 15200 10684 15252 10736
rect 3056 10548 3108 10600
rect 3424 10548 3476 10600
rect 5080 10616 5132 10668
rect 8760 10616 8812 10668
rect 12256 10616 12308 10668
rect 12532 10616 12584 10668
rect 13636 10616 13688 10668
rect 4712 10548 4764 10600
rect 9956 10548 10008 10600
rect 13268 10548 13320 10600
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 14188 10616 14240 10668
rect 15016 10616 15068 10668
rect 14648 10548 14700 10600
rect 14924 10548 14976 10600
rect 15384 10548 15436 10600
rect 4528 10480 4580 10532
rect 4896 10480 4948 10532
rect 5356 10480 5408 10532
rect 12624 10480 12676 10532
rect 17960 10480 18012 10532
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 11796 10412 11848 10464
rect 14004 10412 14056 10464
rect 17776 10412 17828 10464
rect 18420 10455 18472 10464
rect 18420 10421 18429 10455
rect 18429 10421 18463 10455
rect 18463 10421 18472 10455
rect 18420 10412 18472 10421
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 11950 10310 12002 10362
rect 12014 10310 12066 10362
rect 12078 10310 12130 10362
rect 12142 10310 12194 10362
rect 12206 10310 12258 10362
rect 16950 10310 17002 10362
rect 17014 10310 17066 10362
rect 17078 10310 17130 10362
rect 17142 10310 17194 10362
rect 17206 10310 17258 10362
rect 1492 10208 1544 10260
rect 848 10004 900 10056
rect 1768 10004 1820 10056
rect 1584 9936 1636 9988
rect 3700 9868 3752 9920
rect 4068 9868 4120 9920
rect 17776 10251 17828 10260
rect 17776 10217 17785 10251
rect 17785 10217 17819 10251
rect 17819 10217 17828 10251
rect 17776 10208 17828 10217
rect 4988 10140 5040 10192
rect 5080 10183 5132 10192
rect 5080 10149 5089 10183
rect 5089 10149 5123 10183
rect 5123 10149 5132 10183
rect 5080 10140 5132 10149
rect 7564 10072 7616 10124
rect 11152 10140 11204 10192
rect 4988 10004 5040 10056
rect 9772 9936 9824 9988
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 14924 10140 14976 10192
rect 15384 10140 15436 10192
rect 16580 10140 16632 10192
rect 12624 10072 12676 10124
rect 13636 10072 13688 10124
rect 11888 10004 11940 10056
rect 14004 10004 14056 10056
rect 11336 9936 11388 9988
rect 13820 9936 13872 9988
rect 8208 9868 8260 9920
rect 10968 9911 11020 9920
rect 10968 9877 10977 9911
rect 10977 9877 11011 9911
rect 11011 9877 11020 9911
rect 10968 9868 11020 9877
rect 14280 9868 14332 9920
rect 16856 10072 16908 10124
rect 15108 10047 15160 10056
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 15108 10004 15160 10013
rect 15200 10004 15252 10056
rect 17960 10140 18012 10192
rect 17868 10115 17920 10124
rect 17868 10081 17877 10115
rect 17877 10081 17911 10115
rect 17911 10081 17920 10115
rect 17868 10072 17920 10081
rect 15384 9979 15436 9988
rect 15384 9945 15393 9979
rect 15393 9945 15427 9979
rect 15427 9945 15436 9979
rect 15384 9936 15436 9945
rect 16396 9979 16448 9988
rect 16396 9945 16405 9979
rect 16405 9945 16439 9979
rect 16439 9945 16448 9979
rect 16396 9936 16448 9945
rect 17040 9936 17092 9988
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 18420 9868 18472 9920
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 17610 9766 17662 9818
rect 17674 9766 17726 9818
rect 17738 9766 17790 9818
rect 17802 9766 17854 9818
rect 17866 9766 17918 9818
rect 3148 9664 3200 9716
rect 5356 9707 5408 9716
rect 5356 9673 5381 9707
rect 5381 9673 5408 9707
rect 5356 9664 5408 9673
rect 7288 9664 7340 9716
rect 8300 9664 8352 9716
rect 9956 9664 10008 9716
rect 11888 9664 11940 9716
rect 13728 9664 13780 9716
rect 15384 9664 15436 9716
rect 16028 9664 16080 9716
rect 3056 9596 3108 9648
rect 5264 9596 5316 9648
rect 848 9528 900 9580
rect 2228 9528 2280 9580
rect 2872 9528 2924 9580
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 4528 9460 4580 9512
rect 10048 9596 10100 9648
rect 16580 9664 16632 9716
rect 16764 9664 16816 9716
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 6092 9528 6144 9580
rect 6644 9528 6696 9580
rect 6920 9528 6972 9580
rect 9680 9528 9732 9580
rect 10784 9528 10836 9580
rect 15200 9528 15252 9580
rect 15384 9528 15436 9580
rect 15752 9528 15804 9580
rect 5724 9503 5776 9512
rect 5724 9469 5733 9503
rect 5733 9469 5767 9503
rect 5767 9469 5776 9503
rect 5724 9460 5776 9469
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 5908 9503 5960 9512
rect 5908 9469 5917 9503
rect 5917 9469 5951 9503
rect 5951 9469 5960 9503
rect 5908 9460 5960 9469
rect 6460 9460 6512 9512
rect 1860 9324 1912 9376
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 3608 9392 3660 9444
rect 3976 9392 4028 9444
rect 5080 9324 5132 9376
rect 5632 9392 5684 9444
rect 6644 9392 6696 9444
rect 9036 9460 9088 9512
rect 16580 9528 16632 9580
rect 16948 9528 17000 9580
rect 18328 9571 18380 9580
rect 18328 9537 18337 9571
rect 18337 9537 18371 9571
rect 18371 9537 18380 9571
rect 18328 9528 18380 9537
rect 10416 9392 10468 9444
rect 15016 9392 15068 9444
rect 15936 9324 15988 9376
rect 16304 9324 16356 9376
rect 17132 9460 17184 9512
rect 17868 9460 17920 9512
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 18420 9392 18472 9444
rect 17592 9324 17644 9376
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 11950 9222 12002 9274
rect 12014 9222 12066 9274
rect 12078 9222 12130 9274
rect 12142 9222 12194 9274
rect 12206 9222 12258 9274
rect 16950 9222 17002 9274
rect 17014 9222 17066 9274
rect 17078 9222 17130 9274
rect 17142 9222 17194 9274
rect 17206 9222 17258 9274
rect 5540 9120 5592 9172
rect 5816 9120 5868 9172
rect 13084 9120 13136 9172
rect 13268 9120 13320 9172
rect 15108 9120 15160 9172
rect 18052 9120 18104 9172
rect 4160 9052 4212 9104
rect 15752 9052 15804 9104
rect 3148 8984 3200 9036
rect 3516 8984 3568 9036
rect 4988 8984 5040 9036
rect 6644 8984 6696 9036
rect 1492 8916 1544 8968
rect 1676 8916 1728 8968
rect 2872 8916 2924 8968
rect 8576 8916 8628 8968
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 11704 8984 11756 9036
rect 12348 8984 12400 9036
rect 14188 8984 14240 9036
rect 15384 8984 15436 9036
rect 17500 8984 17552 9036
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 3148 8848 3200 8900
rect 7288 8848 7340 8900
rect 8392 8848 8444 8900
rect 15200 8916 15252 8968
rect 17960 8959 18012 8968
rect 17960 8925 17969 8959
rect 17969 8925 18003 8959
rect 18003 8925 18012 8959
rect 17960 8916 18012 8925
rect 18880 8984 18932 9036
rect 17500 8848 17552 8900
rect 7012 8780 7064 8832
rect 14648 8780 14700 8832
rect 15016 8780 15068 8832
rect 17592 8780 17644 8832
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 17610 8678 17662 8730
rect 17674 8678 17726 8730
rect 17738 8678 17790 8730
rect 17802 8678 17854 8730
rect 17866 8678 17918 8730
rect 4160 8619 4212 8628
rect 4160 8585 4169 8619
rect 4169 8585 4203 8619
rect 4203 8585 4212 8619
rect 4160 8576 4212 8585
rect 5724 8576 5776 8628
rect 7380 8576 7432 8628
rect 7932 8576 7984 8628
rect 8484 8576 8536 8628
rect 4804 8508 4856 8560
rect 6644 8551 6696 8560
rect 6644 8517 6653 8551
rect 6653 8517 6687 8551
rect 6687 8517 6696 8551
rect 6644 8508 6696 8517
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 4068 8440 4120 8492
rect 5172 8440 5224 8492
rect 6092 8440 6144 8492
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 9588 8508 9640 8560
rect 11152 8576 11204 8628
rect 11336 8576 11388 8628
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 14372 8576 14424 8628
rect 18052 8576 18104 8628
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 3056 8372 3108 8424
rect 4804 8372 4856 8424
rect 4988 8372 5040 8424
rect 6644 8372 6696 8424
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 7656 8440 7708 8492
rect 10048 8440 10100 8492
rect 10876 8440 10928 8492
rect 11520 8440 11572 8492
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13728 8372 13780 8424
rect 14832 8440 14884 8492
rect 15660 8440 15712 8492
rect 14464 8372 14516 8424
rect 14740 8372 14792 8424
rect 4436 8279 4488 8288
rect 4436 8245 4445 8279
rect 4445 8245 4479 8279
rect 4479 8245 4488 8279
rect 4436 8236 4488 8245
rect 6460 8236 6512 8288
rect 7196 8236 7248 8288
rect 7564 8304 7616 8356
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 8944 8304 8996 8356
rect 9680 8347 9732 8356
rect 9680 8313 9689 8347
rect 9689 8313 9723 8347
rect 9723 8313 9732 8347
rect 9680 8304 9732 8313
rect 10508 8304 10560 8356
rect 7472 8236 7524 8245
rect 9772 8236 9824 8288
rect 12532 8236 12584 8288
rect 14464 8236 14516 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 11950 8134 12002 8186
rect 12014 8134 12066 8186
rect 12078 8134 12130 8186
rect 12142 8134 12194 8186
rect 12206 8134 12258 8186
rect 16950 8134 17002 8186
rect 17014 8134 17066 8186
rect 17078 8134 17130 8186
rect 17142 8134 17194 8186
rect 17206 8134 17258 8186
rect 2412 8032 2464 8084
rect 5908 8032 5960 8084
rect 7196 8032 7248 8084
rect 7656 8032 7708 8084
rect 11520 8032 11572 8084
rect 17500 8032 17552 8084
rect 3976 7964 4028 8016
rect 3608 7896 3660 7948
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 2504 7828 2556 7880
rect 2964 7828 3016 7880
rect 4160 7828 4212 7880
rect 4252 7760 4304 7812
rect 1584 7692 1636 7744
rect 3424 7692 3476 7744
rect 16304 7964 16356 8016
rect 4804 7896 4856 7948
rect 7104 7896 7156 7948
rect 7748 7828 7800 7880
rect 8484 7896 8536 7948
rect 10140 7896 10192 7948
rect 14188 7896 14240 7948
rect 8208 7828 8260 7880
rect 8576 7828 8628 7880
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 9220 7760 9272 7812
rect 6368 7692 6420 7744
rect 6644 7692 6696 7744
rect 7564 7692 7616 7744
rect 8300 7692 8352 7744
rect 13636 7692 13688 7744
rect 14832 7692 14884 7744
rect 18972 7692 19024 7744
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 17610 7590 17662 7642
rect 17674 7590 17726 7642
rect 17738 7590 17790 7642
rect 17802 7590 17854 7642
rect 17866 7590 17918 7642
rect 4988 7488 5040 7540
rect 5264 7488 5316 7540
rect 1768 7420 1820 7472
rect 7104 7420 7156 7472
rect 848 7352 900 7404
rect 7840 7352 7892 7404
rect 8484 7488 8536 7540
rect 13912 7488 13964 7540
rect 16856 7488 16908 7540
rect 11152 7420 11204 7472
rect 11428 7420 11480 7472
rect 12440 7420 12492 7472
rect 13636 7420 13688 7472
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 16856 7352 16908 7404
rect 11152 7284 11204 7336
rect 14004 7284 14056 7336
rect 16304 7327 16356 7336
rect 16304 7293 16313 7327
rect 16313 7293 16347 7327
rect 16347 7293 16356 7327
rect 16304 7284 16356 7293
rect 6184 7216 6236 7268
rect 1676 7148 1728 7200
rect 2504 7148 2556 7200
rect 7196 7148 7248 7200
rect 7472 7148 7524 7200
rect 11336 7148 11388 7200
rect 14464 7148 14516 7200
rect 15200 7148 15252 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 11950 7046 12002 7098
rect 12014 7046 12066 7098
rect 12078 7046 12130 7098
rect 12142 7046 12194 7098
rect 12206 7046 12258 7098
rect 16950 7046 17002 7098
rect 17014 7046 17066 7098
rect 17078 7046 17130 7098
rect 17142 7046 17194 7098
rect 17206 7046 17258 7098
rect 6552 6944 6604 6996
rect 6920 6944 6972 6996
rect 7840 6944 7892 6996
rect 9312 6944 9364 6996
rect 4160 6876 4212 6928
rect 7012 6876 7064 6928
rect 10876 6944 10928 6996
rect 16304 6944 16356 6996
rect 2412 6808 2464 6860
rect 8392 6808 8444 6860
rect 10140 6808 10192 6860
rect 12348 6808 12400 6860
rect 1768 6740 1820 6792
rect 3056 6740 3108 6792
rect 4160 6740 4212 6792
rect 4988 6783 5040 6792
rect 4988 6749 4997 6783
rect 4997 6749 5031 6783
rect 5031 6749 5040 6783
rect 4988 6740 5040 6749
rect 9772 6740 9824 6792
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 11060 6740 11112 6792
rect 12532 6783 12584 6792
rect 12532 6749 12541 6783
rect 12541 6749 12575 6783
rect 12575 6749 12584 6783
rect 12532 6740 12584 6749
rect 16028 6876 16080 6928
rect 16120 6876 16172 6928
rect 14004 6808 14056 6860
rect 2964 6715 3016 6724
rect 2964 6681 2973 6715
rect 2973 6681 3007 6715
rect 3007 6681 3016 6715
rect 2964 6672 3016 6681
rect 6828 6672 6880 6724
rect 8944 6672 8996 6724
rect 3332 6604 3384 6656
rect 5172 6604 5224 6656
rect 9772 6604 9824 6656
rect 11152 6672 11204 6724
rect 11520 6672 11572 6724
rect 12348 6672 12400 6724
rect 15660 6672 15712 6724
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 18788 6740 18840 6792
rect 16212 6672 16264 6724
rect 9956 6604 10008 6656
rect 14004 6604 14056 6656
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 17610 6502 17662 6554
rect 17674 6502 17726 6554
rect 17738 6502 17790 6554
rect 17802 6502 17854 6554
rect 17866 6502 17918 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 5816 6400 5868 6452
rect 9680 6400 9732 6452
rect 9772 6400 9824 6452
rect 1400 6375 1452 6384
rect 1400 6341 1409 6375
rect 1409 6341 1443 6375
rect 1443 6341 1452 6375
rect 1400 6332 1452 6341
rect 2320 6332 2372 6384
rect 2964 6332 3016 6384
rect 10140 6332 10192 6384
rect 10600 6400 10652 6452
rect 18144 6400 18196 6452
rect 10692 6332 10744 6384
rect 13728 6375 13780 6384
rect 13728 6341 13737 6375
rect 13737 6341 13771 6375
rect 13771 6341 13780 6375
rect 13728 6332 13780 6341
rect 940 6264 992 6316
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 7012 6307 7064 6316
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 8852 6264 8904 6316
rect 9496 6264 9548 6316
rect 1400 6196 1452 6248
rect 10048 6196 10100 6248
rect 1768 6171 1820 6180
rect 1768 6137 1777 6171
rect 1777 6137 1811 6171
rect 1811 6137 1820 6171
rect 1768 6128 1820 6137
rect 4712 6128 4764 6180
rect 9956 6128 10008 6180
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 6184 6060 6236 6112
rect 10232 6103 10284 6112
rect 10232 6069 10241 6103
rect 10241 6069 10275 6103
rect 10275 6069 10284 6103
rect 14280 6264 14332 6316
rect 16304 6264 16356 6316
rect 16488 6264 16540 6316
rect 11796 6196 11848 6248
rect 12348 6196 12400 6248
rect 10232 6060 10284 6069
rect 10692 6060 10744 6112
rect 12440 6060 12492 6112
rect 13820 6196 13872 6248
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 18236 6239 18288 6248
rect 18236 6205 18245 6239
rect 18245 6205 18279 6239
rect 18279 6205 18288 6239
rect 18236 6196 18288 6205
rect 13360 6171 13412 6180
rect 13360 6137 13369 6171
rect 13369 6137 13403 6171
rect 13403 6137 13412 6171
rect 13360 6128 13412 6137
rect 15844 6171 15896 6180
rect 15844 6137 15853 6171
rect 15853 6137 15887 6171
rect 15887 6137 15896 6171
rect 15844 6128 15896 6137
rect 16212 6128 16264 6180
rect 16488 6128 16540 6180
rect 16764 6128 16816 6180
rect 18328 6060 18380 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 11950 5958 12002 6010
rect 12014 5958 12066 6010
rect 12078 5958 12130 6010
rect 12142 5958 12194 6010
rect 12206 5958 12258 6010
rect 16950 5958 17002 6010
rect 17014 5958 17066 6010
rect 17078 5958 17130 6010
rect 17142 5958 17194 6010
rect 17206 5958 17258 6010
rect 2320 5856 2372 5908
rect 3240 5856 3292 5908
rect 4068 5856 4120 5908
rect 4344 5856 4396 5908
rect 6644 5856 6696 5908
rect 4712 5788 4764 5840
rect 8116 5788 8168 5840
rect 13176 5856 13228 5908
rect 11428 5720 11480 5772
rect 13820 5788 13872 5840
rect 4528 5652 4580 5704
rect 10876 5652 10928 5704
rect 9312 5584 9364 5636
rect 12348 5652 12400 5704
rect 13544 5652 13596 5704
rect 14280 5652 14332 5704
rect 14832 5856 14884 5908
rect 15016 5856 15068 5908
rect 16580 5856 16632 5908
rect 15936 5720 15988 5772
rect 14832 5695 14884 5704
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 15384 5652 15436 5704
rect 16488 5720 16540 5772
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 16488 5584 16540 5636
rect 18236 5584 18288 5636
rect 13544 5516 13596 5568
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 16212 5559 16264 5568
rect 16212 5525 16221 5559
rect 16221 5525 16255 5559
rect 16255 5525 16264 5559
rect 16212 5516 16264 5525
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 17610 5414 17662 5466
rect 17674 5414 17726 5466
rect 17738 5414 17790 5466
rect 17802 5414 17854 5466
rect 17866 5414 17918 5466
rect 1492 5312 1544 5364
rect 4160 5312 4212 5364
rect 7380 5312 7432 5364
rect 8024 5355 8076 5364
rect 8024 5321 8033 5355
rect 8033 5321 8067 5355
rect 8067 5321 8076 5355
rect 8024 5312 8076 5321
rect 11060 5312 11112 5364
rect 10876 5244 10928 5296
rect 848 5176 900 5228
rect 6828 5176 6880 5228
rect 7380 5176 7432 5228
rect 7748 5219 7800 5228
rect 7748 5185 7757 5219
rect 7757 5185 7791 5219
rect 7791 5185 7800 5219
rect 7748 5176 7800 5185
rect 5172 5083 5224 5092
rect 5172 5049 5181 5083
rect 5181 5049 5215 5083
rect 5215 5049 5224 5083
rect 5172 5040 5224 5049
rect 6920 5040 6972 5092
rect 7748 5040 7800 5092
rect 8024 5108 8076 5160
rect 8300 5176 8352 5228
rect 12256 5176 12308 5228
rect 12992 5287 13044 5296
rect 12992 5253 13001 5287
rect 13001 5253 13035 5287
rect 13035 5253 13044 5287
rect 12992 5244 13044 5253
rect 14556 5244 14608 5296
rect 16212 5312 16264 5364
rect 16396 5244 16448 5296
rect 13268 5176 13320 5228
rect 13452 5219 13504 5228
rect 13452 5185 13461 5219
rect 13461 5185 13495 5219
rect 13495 5185 13504 5219
rect 13452 5176 13504 5185
rect 13728 5219 13780 5228
rect 13728 5185 13737 5219
rect 13737 5185 13771 5219
rect 13771 5185 13780 5219
rect 13728 5176 13780 5185
rect 15292 5176 15344 5228
rect 15384 5219 15436 5228
rect 15384 5185 15393 5219
rect 15393 5185 15427 5219
rect 15427 5185 15436 5219
rect 15384 5176 15436 5185
rect 13176 5151 13228 5160
rect 13176 5117 13185 5151
rect 13185 5117 13219 5151
rect 13219 5117 13228 5151
rect 13176 5108 13228 5117
rect 11060 5040 11112 5092
rect 11704 5040 11756 5092
rect 3056 4972 3108 5024
rect 8300 4972 8352 5024
rect 9036 4972 9088 5024
rect 9312 4972 9364 5024
rect 11152 4972 11204 5024
rect 11428 4972 11480 5024
rect 16764 4972 16816 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 11950 4870 12002 4922
rect 12014 4870 12066 4922
rect 12078 4870 12130 4922
rect 12142 4870 12194 4922
rect 12206 4870 12258 4922
rect 16950 4870 17002 4922
rect 17014 4870 17066 4922
rect 17078 4870 17130 4922
rect 17142 4870 17194 4922
rect 17206 4870 17258 4922
rect 1492 4700 1544 4752
rect 13728 4768 13780 4820
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 4068 4700 4120 4752
rect 12072 4743 12124 4752
rect 12072 4709 12081 4743
rect 12081 4709 12115 4743
rect 12115 4709 12124 4743
rect 12072 4700 12124 4709
rect 12440 4743 12492 4752
rect 12440 4709 12449 4743
rect 12449 4709 12483 4743
rect 12483 4709 12492 4743
rect 12440 4700 12492 4709
rect 13084 4700 13136 4752
rect 6828 4632 6880 4684
rect 8944 4632 8996 4684
rect 9220 4675 9272 4684
rect 9220 4641 9229 4675
rect 9229 4641 9263 4675
rect 9263 4641 9272 4675
rect 9220 4632 9272 4641
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 10232 4632 10284 4684
rect 12532 4675 12584 4684
rect 12532 4641 12541 4675
rect 12541 4641 12575 4675
rect 12575 4641 12584 4675
rect 12532 4632 12584 4641
rect 13820 4632 13872 4684
rect 16304 4768 16356 4820
rect 16672 4811 16724 4820
rect 16672 4777 16681 4811
rect 16681 4777 16715 4811
rect 16715 4777 16724 4811
rect 16672 4768 16724 4777
rect 16856 4768 16908 4820
rect 8852 4564 8904 4616
rect 7748 4496 7800 4548
rect 9036 4496 9088 4548
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 11612 4564 11664 4616
rect 14464 4564 14516 4616
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 18512 4700 18564 4752
rect 15660 4564 15712 4573
rect 11152 4496 11204 4548
rect 8944 4471 8996 4480
rect 8944 4437 8953 4471
rect 8953 4437 8987 4471
rect 8987 4437 8996 4471
rect 8944 4428 8996 4437
rect 9312 4428 9364 4480
rect 12348 4496 12400 4548
rect 16764 4607 16816 4616
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 16304 4539 16356 4548
rect 16304 4505 16313 4539
rect 16313 4505 16347 4539
rect 16347 4505 16356 4539
rect 16304 4496 16356 4505
rect 16396 4539 16448 4548
rect 16396 4505 16405 4539
rect 16405 4505 16439 4539
rect 16439 4505 16448 4539
rect 16396 4496 16448 4505
rect 13820 4428 13872 4480
rect 14004 4428 14056 4480
rect 14924 4428 14976 4480
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 17610 4326 17662 4378
rect 17674 4326 17726 4378
rect 17738 4326 17790 4378
rect 17802 4326 17854 4378
rect 17866 4326 17918 4378
rect 2412 4224 2464 4276
rect 9312 4224 9364 4276
rect 9864 4224 9916 4276
rect 10140 4267 10192 4276
rect 10140 4233 10149 4267
rect 10149 4233 10183 4267
rect 10183 4233 10192 4267
rect 10140 4224 10192 4233
rect 3148 4199 3200 4208
rect 3148 4165 3157 4199
rect 3157 4165 3191 4199
rect 3191 4165 3200 4199
rect 3148 4156 3200 4165
rect 9956 4156 10008 4208
rect 11060 4156 11112 4208
rect 14740 4199 14792 4208
rect 14740 4165 14749 4199
rect 14749 4165 14783 4199
rect 14783 4165 14792 4199
rect 14740 4156 14792 4165
rect 15108 4156 15160 4208
rect 16396 4156 16448 4208
rect 17500 4199 17552 4208
rect 17500 4165 17509 4199
rect 17509 4165 17543 4199
rect 17543 4165 17552 4199
rect 17500 4156 17552 4165
rect 17960 4156 18012 4208
rect 848 4088 900 4140
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 8760 4088 8812 4140
rect 10140 4088 10192 4140
rect 15200 4088 15252 4140
rect 15292 4088 15344 4140
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 18328 4020 18380 4072
rect 1860 3952 1912 4004
rect 5816 3995 5868 4004
rect 5816 3961 5825 3995
rect 5825 3961 5859 3995
rect 5859 3961 5868 3995
rect 5816 3952 5868 3961
rect 10324 3952 10376 4004
rect 12348 3952 12400 4004
rect 3240 3884 3292 3936
rect 9404 3884 9456 3936
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 16212 3884 16264 3936
rect 18420 3927 18472 3936
rect 18420 3893 18429 3927
rect 18429 3893 18463 3927
rect 18463 3893 18472 3927
rect 18420 3884 18472 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 11950 3782 12002 3834
rect 12014 3782 12066 3834
rect 12078 3782 12130 3834
rect 12142 3782 12194 3834
rect 12206 3782 12258 3834
rect 16950 3782 17002 3834
rect 17014 3782 17066 3834
rect 17078 3782 17130 3834
rect 17142 3782 17194 3834
rect 17206 3782 17258 3834
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 7288 3680 7340 3732
rect 5080 3612 5132 3664
rect 1860 3544 1912 3596
rect 15108 3680 15160 3732
rect 17316 3680 17368 3732
rect 3608 3476 3660 3528
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 4252 3408 4304 3460
rect 13452 3612 13504 3664
rect 11152 3544 11204 3596
rect 14464 3544 14516 3596
rect 15476 3544 15528 3596
rect 9588 3476 9640 3528
rect 11336 3476 11388 3528
rect 12164 3476 12216 3528
rect 13084 3476 13136 3528
rect 11244 3408 11296 3460
rect 10968 3340 11020 3392
rect 12532 3340 12584 3392
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 17610 3238 17662 3290
rect 17674 3238 17726 3290
rect 17738 3238 17790 3290
rect 17802 3238 17854 3290
rect 17866 3238 17918 3290
rect 1676 3111 1728 3120
rect 1676 3077 1685 3111
rect 1685 3077 1719 3111
rect 1719 3077 1728 3111
rect 1676 3068 1728 3077
rect 848 3000 900 3052
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 9588 3136 9640 3188
rect 10968 3136 11020 3188
rect 3976 3068 4028 3120
rect 4252 3068 4304 3120
rect 6460 3068 6512 3120
rect 4804 3000 4856 3052
rect 8852 3000 8904 3052
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 10508 3000 10560 3052
rect 10692 3000 10744 3052
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11428 3000 11480 3052
rect 12348 3111 12400 3120
rect 12348 3077 12357 3111
rect 12357 3077 12391 3111
rect 12391 3077 12400 3111
rect 12348 3068 12400 3077
rect 13912 3068 13964 3120
rect 15016 3068 15068 3120
rect 12164 3043 12216 3052
rect 12164 3009 12171 3043
rect 12171 3009 12216 3043
rect 12164 3000 12216 3009
rect 12532 3000 12584 3052
rect 14556 3043 14608 3052
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 7380 2864 7432 2916
rect 14648 2932 14700 2984
rect 2320 2839 2372 2848
rect 2320 2805 2329 2839
rect 2329 2805 2363 2839
rect 2363 2805 2372 2839
rect 2320 2796 2372 2805
rect 8208 2796 8260 2848
rect 18696 2796 18748 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 11950 2694 12002 2746
rect 12014 2694 12066 2746
rect 12078 2694 12130 2746
rect 12142 2694 12194 2746
rect 12206 2694 12258 2746
rect 16950 2694 17002 2746
rect 17014 2694 17066 2746
rect 17078 2694 17130 2746
rect 17142 2694 17194 2746
rect 17206 2694 17258 2746
rect 4620 2592 4672 2644
rect 11060 2592 11112 2644
rect 15568 2592 15620 2644
rect 1308 2524 1360 2576
rect 10784 2524 10836 2576
rect 15292 2524 15344 2576
rect 17408 2524 17460 2576
rect 10692 2456 10744 2508
rect 17500 2456 17552 2508
rect 1216 2320 1268 2372
rect 7472 2388 7524 2440
rect 8944 2431 8996 2440
rect 8944 2397 8953 2431
rect 8953 2397 8987 2431
rect 8987 2397 8996 2431
rect 8944 2388 8996 2397
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16580 2388 16632 2440
rect 18604 2388 18656 2440
rect 3332 2320 3384 2372
rect 9956 2320 10008 2372
rect 13728 2320 13780 2372
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 16212 2320 16264 2372
rect 18052 2363 18104 2372
rect 18052 2329 18061 2363
rect 18061 2329 18095 2363
rect 18095 2329 18104 2363
rect 18052 2320 18104 2329
rect 18420 2295 18472 2304
rect 18420 2261 18429 2295
rect 18429 2261 18463 2295
rect 18463 2261 18472 2295
rect 18420 2252 18472 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 17610 2150 17662 2202
rect 17674 2150 17726 2202
rect 17738 2150 17790 2202
rect 17802 2150 17854 2202
rect 17866 2150 17918 2202
<< metal2 >>
rect 17866 18592 17922 18601
rect 17866 18527 17922 18536
rect 1858 18048 1914 18057
rect 1858 17983 1914 17992
rect 1872 17270 1900 17983
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 17880 17626 17908 18527
rect 18144 17672 18196 17678
rect 2610 17436 2918 17445
rect 2610 17434 2616 17436
rect 2672 17434 2696 17436
rect 2752 17434 2776 17436
rect 2832 17434 2856 17436
rect 2912 17434 2918 17436
rect 2672 17382 2674 17434
rect 2854 17382 2856 17434
rect 2610 17380 2616 17382
rect 2672 17380 2696 17382
rect 2752 17380 2776 17382
rect 2832 17380 2856 17382
rect 2912 17380 2918 17382
rect 2610 17371 2918 17380
rect 1860 17264 1912 17270
rect 1860 17206 1912 17212
rect 848 17196 900 17202
rect 848 17138 900 17144
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 860 17105 888 17138
rect 846 17096 902 17105
rect 846 17031 902 17040
rect 2320 17060 2372 17066
rect 2320 17002 2372 17008
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1032 16176 1084 16182
rect 1032 16118 1084 16124
rect 1044 15881 1072 16118
rect 1030 15872 1086 15881
rect 1412 15858 1440 16934
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1490 16008 1546 16017
rect 1490 15943 1492 15952
rect 1544 15943 1546 15952
rect 1492 15914 1544 15920
rect 1412 15830 1532 15858
rect 1030 15807 1086 15816
rect 848 15020 900 15026
rect 848 14962 900 14968
rect 860 14929 888 14962
rect 846 14920 902 14929
rect 846 14855 902 14864
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1504 13546 1532 15830
rect 1412 13518 1532 13546
rect 848 12844 900 12850
rect 848 12786 900 12792
rect 860 12753 888 12786
rect 846 12744 902 12753
rect 846 12679 902 12688
rect 848 11756 900 11762
rect 848 11698 900 11704
rect 860 11665 888 11698
rect 846 11656 902 11665
rect 846 11591 902 11600
rect 1306 11248 1362 11257
rect 1306 11183 1362 11192
rect 1214 10704 1270 10713
rect 1214 10639 1270 10648
rect 846 10296 902 10305
rect 846 10231 902 10240
rect 860 10062 888 10231
rect 848 10056 900 10062
rect 848 9998 900 10004
rect 848 9580 900 9586
rect 848 9522 900 9528
rect 860 9489 888 9522
rect 846 9480 902 9489
rect 846 9415 902 9424
rect 848 7404 900 7410
rect 848 7346 900 7352
rect 860 7313 888 7346
rect 846 7304 902 7313
rect 846 7239 902 7248
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 952 6089 980 6258
rect 938 6080 994 6089
rect 938 6015 994 6024
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5137 888 5170
rect 846 5128 902 5137
rect 846 5063 902 5072
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 860 4049 888 4082
rect 846 4040 902 4049
rect 846 3975 902 3984
rect 848 3052 900 3058
rect 848 2994 900 3000
rect 860 2961 888 2994
rect 846 2952 902 2961
rect 846 2887 902 2896
rect 1228 2378 1256 10639
rect 1320 2582 1348 11183
rect 1412 10033 1440 13518
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1504 11558 1532 12922
rect 1596 12442 1624 16050
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1492 11280 1544 11286
rect 1492 11222 1544 11228
rect 1504 10554 1532 11222
rect 1596 10742 1624 12378
rect 1688 11286 1716 13738
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1780 12374 1808 13670
rect 1872 12986 1900 14554
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 1768 12368 1820 12374
rect 1768 12310 1820 12316
rect 1676 11280 1728 11286
rect 1676 11222 1728 11228
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1584 10736 1636 10742
rect 1584 10678 1636 10684
rect 1688 10674 1716 11086
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1504 10526 1624 10554
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1504 10266 1532 10406
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1398 10024 1454 10033
rect 1596 9994 1624 10526
rect 1398 9959 1454 9968
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1504 8106 1532 8910
rect 1412 8078 1532 8106
rect 1412 6390 1440 8078
rect 1596 7834 1624 9930
rect 1688 8974 1716 10610
rect 1780 10062 1808 12310
rect 2332 12238 2360 17002
rect 2516 16114 2544 17138
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 4172 16726 4200 17002
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 2610 16348 2918 16357
rect 2610 16346 2616 16348
rect 2672 16346 2696 16348
rect 2752 16346 2776 16348
rect 2832 16346 2856 16348
rect 2912 16346 2918 16348
rect 2672 16294 2674 16346
rect 2854 16294 2856 16346
rect 2610 16292 2616 16294
rect 2672 16292 2696 16294
rect 2752 16292 2776 16294
rect 2832 16292 2856 16294
rect 2912 16292 2918 16294
rect 2610 16283 2918 16292
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1872 10674 1900 12038
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1964 10554 1992 10610
rect 1872 10526 1992 10554
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1872 9466 1900 10526
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 2228 9580 2280 9586
rect 2332 9568 2360 11494
rect 2280 9540 2360 9568
rect 2228 9522 2280 9528
rect 1780 9438 1900 9466
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1504 7806 1624 7834
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 1412 6254 1440 6326
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1504 5370 1532 7806
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 6118 1624 7686
rect 1780 7478 1808 9438
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1768 7472 1820 7478
rect 1768 7414 1820 7420
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1504 4758 1532 5306
rect 1492 4752 1544 4758
rect 1492 4694 1544 4700
rect 1688 3126 1716 7142
rect 1780 6798 1808 7414
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1766 6216 1822 6225
rect 1766 6151 1768 6160
rect 1820 6151 1822 6160
rect 1768 6122 1820 6128
rect 1872 4010 1900 9318
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2332 7970 2360 9540
rect 2424 8090 2452 15506
rect 2976 15434 3004 16186
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3068 16017 3096 16050
rect 3054 16008 3110 16017
rect 3054 15943 3110 15952
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 2976 13326 3004 15370
rect 2964 13320 3016 13326
rect 3016 13280 3096 13308
rect 2964 13262 3016 13268
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 2502 10024 2558 10033
rect 2502 9959 2558 9968
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2516 7970 2544 9959
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 8945 2636 9318
rect 2884 8974 2912 9522
rect 2872 8968 2924 8974
rect 2594 8936 2650 8945
rect 2872 8910 2924 8916
rect 2594 8871 2650 8880
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2240 7942 2360 7970
rect 2424 7942 2544 7970
rect 2240 7698 2268 7942
rect 2320 7880 2372 7886
rect 2318 7848 2320 7857
rect 2372 7848 2374 7857
rect 2318 7783 2374 7792
rect 2240 7670 2360 7698
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2042 6760 2098 6769
rect 2332 6746 2360 7670
rect 2424 6866 2452 7942
rect 2976 7886 3004 11562
rect 3068 10606 3096 13280
rect 3160 12434 3188 16050
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3436 13870 3464 14758
rect 3424 13864 3476 13870
rect 3528 13841 3556 14962
rect 3424 13806 3476 13812
rect 3514 13832 3570 13841
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12434 3372 13262
rect 3436 12850 3464 13806
rect 3514 13767 3570 13776
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3160 12406 3280 12434
rect 3344 12406 3556 12434
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3146 9752 3202 9761
rect 3146 9687 3148 9696
rect 3200 9687 3202 9696
rect 3148 9658 3200 9664
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3068 8430 3096 9590
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3160 9042 3188 9522
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2516 7206 2544 7822
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 3068 6798 3096 8366
rect 3056 6792 3108 6798
rect 2332 6718 2452 6746
rect 3056 6734 3108 6740
rect 2042 6695 2098 6704
rect 2056 6458 2084 6695
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2332 5914 2360 6326
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2424 4282 2452 6718
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2976 6390 3004 6666
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 3068 5030 3096 6734
rect 3160 5794 3188 8842
rect 3252 5914 3280 12406
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3344 11354 3372 12174
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3344 9586 3372 11290
rect 3528 10674 3556 12406
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3344 6662 3372 9522
rect 3436 8401 3464 10542
rect 3528 9042 3556 10610
rect 3620 9450 3648 13194
rect 3712 9926 3740 16458
rect 4710 16416 4766 16425
rect 4710 16351 4766 16360
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3804 12850 3832 13330
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3804 11286 3832 11766
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3790 10840 3846 10849
rect 3790 10775 3846 10784
rect 3804 10742 3832 10775
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3698 9480 3754 9489
rect 3608 9444 3660 9450
rect 3698 9415 3754 9424
rect 3608 9386 3660 9392
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3712 8498 3740 9415
rect 3896 8498 3924 15098
rect 3974 15056 4030 15065
rect 3974 14991 4030 15000
rect 3988 13258 4016 14991
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 4080 11694 4108 16118
rect 4342 15600 4398 15609
rect 4342 15535 4398 15544
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4068 11688 4120 11694
rect 3974 11656 4030 11665
rect 4068 11630 4120 11636
rect 3974 11591 4030 11600
rect 3988 11558 4016 11591
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10810 4016 10950
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3976 10668 4028 10674
rect 4080 10656 4108 11630
rect 4172 10810 4200 14486
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4028 10628 4108 10656
rect 3976 10610 4028 10616
rect 3988 9450 4016 10610
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3422 8392 3478 8401
rect 3422 8327 3478 8336
rect 3436 7750 3464 8327
rect 3620 7954 3648 8434
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3160 5766 3280 5794
rect 3146 5264 3202 5273
rect 3146 5199 3202 5208
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 3160 4214 3188 5199
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1872 3602 1900 3946
rect 3252 3942 3280 5766
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 3620 3534 3648 7890
rect 3896 3738 3924 8434
rect 3988 8022 4016 9386
rect 4080 8945 4108 9862
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4066 8936 4122 8945
rect 4066 8871 4122 8880
rect 4066 8800 4122 8809
rect 4066 8735 4122 8744
rect 4080 8498 4108 8735
rect 4172 8634 4200 9046
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4172 6934 4200 7822
rect 4264 7818 4292 11834
rect 4356 11082 4384 15535
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4434 12880 4490 12889
rect 4540 12850 4568 13126
rect 4434 12815 4436 12824
rect 4488 12815 4490 12824
rect 4528 12844 4580 12850
rect 4436 12786 4488 12792
rect 4528 12786 4580 12792
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4080 4758 4108 5850
rect 4172 5370 4200 6734
rect 4356 5914 4384 11018
rect 4448 8294 4476 11086
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4540 10538 4568 10746
rect 4632 10742 4660 12106
rect 4724 11218 4752 16351
rect 4804 16040 4856 16046
rect 4802 16008 4804 16017
rect 4856 16008 4858 16017
rect 4802 15943 4858 15952
rect 4894 13424 4950 13433
rect 4894 13359 4950 13368
rect 4908 12850 4936 13359
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4540 5710 4568 9454
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 4172 3210 4200 5306
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 3988 3182 4200 3210
rect 3988 3126 4016 3182
rect 4264 3126 4292 3402
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1308 2576 1360 2582
rect 1308 2518 1360 2524
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 1872 1737 1900 2994
rect 2318 2952 2374 2961
rect 2318 2887 2374 2896
rect 2332 2854 2360 2887
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 4632 2650 4660 10678
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4724 6186 4752 10542
rect 4816 8566 4844 11086
rect 5000 10810 5028 16730
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5092 10674 5120 17138
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 13938 5304 16934
rect 5460 16794 5488 17614
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 16580 17604 16632 17610
rect 17880 17598 18000 17626
rect 18144 17614 18196 17620
rect 16580 17546 16632 17552
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 7610 17436 7918 17445
rect 7610 17434 7616 17436
rect 7672 17434 7696 17436
rect 7752 17434 7776 17436
rect 7832 17434 7856 17436
rect 7912 17434 7918 17436
rect 7672 17382 7674 17434
rect 7854 17382 7856 17434
rect 7610 17380 7616 17382
rect 7672 17380 7696 17382
rect 7752 17380 7776 17382
rect 7832 17380 7856 17382
rect 7912 17380 7918 17382
rect 7610 17371 7918 17380
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5552 16590 5580 16934
rect 6950 16892 7258 16901
rect 6950 16890 6956 16892
rect 7012 16890 7036 16892
rect 7092 16890 7116 16892
rect 7172 16890 7196 16892
rect 7252 16890 7258 16892
rect 7012 16838 7014 16890
rect 7194 16838 7196 16890
rect 6950 16836 6956 16838
rect 7012 16836 7036 16838
rect 7092 16836 7116 16838
rect 7172 16836 7196 16838
rect 7252 16836 7258 16838
rect 6950 16827 7258 16836
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 6552 16720 6604 16726
rect 6552 16662 6604 16668
rect 8312 16674 8340 16730
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5354 16008 5410 16017
rect 5354 15943 5410 15952
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5368 11393 5396 15943
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5552 13462 5580 15030
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5644 13308 5672 16186
rect 5724 15632 5776 15638
rect 5724 15574 5776 15580
rect 5736 13326 5764 15574
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 5552 13280 5672 13308
rect 5724 13320 5776 13326
rect 5354 11384 5410 11393
rect 5354 11319 5410 11328
rect 5552 11286 5580 13280
rect 5724 13262 5776 13268
rect 5736 12850 5764 13262
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5368 10810 5396 11018
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5080 10668 5132 10674
rect 5132 10628 5304 10656
rect 5080 10610 5132 10616
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4908 10180 4936 10474
rect 4988 10192 5040 10198
rect 4908 10152 4988 10180
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4816 7954 4844 8366
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4724 5846 4752 6122
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4816 3058 4844 7890
rect 4908 6769 4936 10152
rect 5080 10192 5132 10198
rect 4988 10134 5040 10140
rect 5078 10160 5080 10169
rect 5132 10160 5134 10169
rect 5078 10095 5134 10104
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9042 5028 9998
rect 5276 9654 5304 10628
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5368 9722 5396 10474
rect 5538 10024 5594 10033
rect 5538 9959 5594 9968
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5000 8430 5028 8978
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 5000 6798 5028 7482
rect 4988 6792 5040 6798
rect 4894 6760 4950 6769
rect 4988 6734 5040 6740
rect 4894 6695 4950 6704
rect 5092 3670 5120 9318
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5184 6662 5212 8434
rect 5276 7546 5304 9590
rect 5552 9178 5580 9959
rect 5644 9450 5672 12786
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5736 11150 5764 12650
rect 5828 11762 5856 15302
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5920 12986 5948 14282
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5920 11762 5948 12922
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5828 11558 5856 11698
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5920 11354 5948 11698
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 6012 9586 6040 12038
rect 6104 11014 6132 14758
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6196 12434 6224 13806
rect 6196 12406 6316 12434
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6104 10577 6132 10950
rect 6090 10568 6146 10577
rect 6090 10503 6146 10512
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5736 8634 5764 9454
rect 5828 9178 5856 9454
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5920 8090 5948 9454
rect 6104 8498 6132 9522
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 6196 7274 6224 11766
rect 6184 7268 6236 7274
rect 6184 7210 6236 7216
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5170 5128 5226 5137
rect 5170 5063 5172 5072
rect 5224 5063 5226 5072
rect 5172 5034 5224 5040
rect 5828 4146 5856 6394
rect 6196 6118 6224 7210
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6288 4185 6316 12406
rect 6380 7750 6408 15302
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6472 12238 6500 13670
rect 6564 12434 6592 16662
rect 6828 16652 6880 16658
rect 8312 16646 8616 16674
rect 6828 16594 6880 16600
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6840 16538 6868 16594
rect 8392 16584 8444 16590
rect 6918 16552 6974 16561
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6656 15337 6684 15438
rect 6642 15328 6698 15337
rect 6642 15263 6698 15272
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6656 13530 6684 14962
rect 6748 14890 6776 16526
rect 6840 16510 6918 16538
rect 6840 15586 6868 16510
rect 8392 16526 8444 16532
rect 6918 16487 6974 16496
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7484 16476 8064 16504
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 6950 15804 7258 15813
rect 6950 15802 6956 15804
rect 7012 15802 7036 15804
rect 7092 15802 7116 15804
rect 7172 15802 7196 15804
rect 7252 15802 7258 15804
rect 7012 15750 7014 15802
rect 7194 15750 7196 15802
rect 6950 15748 6956 15750
rect 7012 15748 7036 15750
rect 7092 15748 7116 15750
rect 7172 15748 7196 15750
rect 7252 15748 7258 15750
rect 6950 15739 7258 15748
rect 6840 15558 6960 15586
rect 6932 14906 6960 15558
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6840 14878 6960 14906
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6564 12406 6684 12434
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6472 11354 6500 11698
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6458 11112 6514 11121
rect 6458 11047 6514 11056
rect 6472 11014 6500 11047
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6472 8809 6500 9454
rect 6564 9081 6592 11494
rect 6656 9586 6684 12406
rect 6748 12374 6776 14826
rect 6840 14600 6868 14878
rect 6950 14716 7258 14725
rect 6950 14714 6956 14716
rect 7012 14714 7036 14716
rect 7092 14714 7116 14716
rect 7172 14714 7196 14716
rect 7252 14714 7258 14716
rect 7012 14662 7014 14714
rect 7194 14662 7196 14714
rect 6950 14660 6956 14662
rect 7012 14660 7036 14662
rect 7092 14660 7116 14662
rect 7172 14660 7196 14662
rect 7252 14660 7258 14662
rect 6950 14651 7258 14660
rect 6840 14572 6960 14600
rect 6826 14512 6882 14521
rect 6826 14447 6882 14456
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6734 11384 6790 11393
rect 6734 11319 6790 11328
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6550 9072 6606 9081
rect 6656 9042 6684 9386
rect 6550 9007 6606 9016
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6458 8800 6514 8809
rect 6458 8735 6514 8744
rect 6656 8566 6684 8978
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 6322 6408 7686
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6274 4176 6330 4185
rect 5816 4140 5868 4146
rect 6274 4111 6330 4120
rect 5816 4082 5868 4088
rect 5814 4040 5870 4049
rect 5814 3975 5816 3984
rect 5868 3975 5870 3984
rect 5816 3946 5868 3952
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 6472 3126 6500 8230
rect 6564 7002 6592 8434
rect 6644 8424 6696 8430
rect 6642 8392 6644 8401
rect 6696 8392 6698 8401
rect 6642 8327 6698 8336
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6656 5914 6684 7686
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6748 5817 6776 11319
rect 6840 6730 6868 14447
rect 6932 13802 6960 14572
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 6950 13628 7258 13637
rect 6950 13626 6956 13628
rect 7012 13626 7036 13628
rect 7092 13626 7116 13628
rect 7172 13626 7196 13628
rect 7252 13626 7258 13628
rect 7012 13574 7014 13626
rect 7194 13574 7196 13626
rect 6950 13572 6956 13574
rect 7012 13572 7036 13574
rect 7092 13572 7116 13574
rect 7172 13572 7196 13574
rect 7252 13572 7258 13574
rect 6950 13563 7258 13572
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7024 12753 7052 12786
rect 7208 12753 7236 13466
rect 7010 12744 7066 12753
rect 7010 12679 7066 12688
rect 7194 12744 7250 12753
rect 7300 12714 7328 16390
rect 7194 12679 7250 12688
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 7392 12646 7420 16458
rect 7484 16425 7512 16476
rect 8036 16425 8064 16476
rect 7470 16416 7526 16425
rect 7470 16351 7526 16360
rect 8022 16416 8078 16425
rect 7610 16348 7918 16357
rect 8022 16351 8078 16360
rect 7610 16346 7616 16348
rect 7672 16346 7696 16348
rect 7752 16346 7776 16348
rect 7832 16346 7856 16348
rect 7912 16346 7918 16348
rect 7672 16294 7674 16346
rect 7854 16294 7856 16346
rect 7610 16292 7616 16294
rect 7672 16292 7696 16294
rect 7752 16292 7776 16294
rect 7832 16292 7856 16294
rect 7912 16292 7918 16294
rect 7610 16283 7918 16292
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 7610 15260 7918 15269
rect 7610 15258 7616 15260
rect 7672 15258 7696 15260
rect 7752 15258 7776 15260
rect 7832 15258 7856 15260
rect 7912 15258 7918 15260
rect 7672 15206 7674 15258
rect 7854 15206 7856 15258
rect 7610 15204 7616 15206
rect 7672 15204 7696 15206
rect 7752 15204 7776 15206
rect 7832 15204 7856 15206
rect 7912 15204 7918 15206
rect 7610 15195 7918 15204
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7484 12968 7512 14894
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7576 14482 7604 14758
rect 7668 14618 7696 14962
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 8036 14278 8064 14826
rect 8128 14414 8156 15302
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 7610 14172 7918 14181
rect 7610 14170 7616 14172
rect 7672 14170 7696 14172
rect 7752 14170 7776 14172
rect 7832 14170 7856 14172
rect 7912 14170 7918 14172
rect 7672 14118 7674 14170
rect 7854 14118 7856 14170
rect 7610 14116 7616 14118
rect 7672 14116 7696 14118
rect 7752 14116 7776 14118
rect 7832 14116 7856 14118
rect 7912 14116 7918 14118
rect 7610 14107 7918 14116
rect 8036 14090 8064 14214
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7944 14062 8064 14090
rect 7576 13297 7604 14010
rect 7944 13530 7972 14062
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7562 13288 7618 13297
rect 7562 13223 7618 13232
rect 7610 13084 7918 13093
rect 7610 13082 7616 13084
rect 7672 13082 7696 13084
rect 7752 13082 7776 13084
rect 7832 13082 7856 13084
rect 7912 13082 7918 13084
rect 7672 13030 7674 13082
rect 7854 13030 7856 13082
rect 7610 13028 7616 13030
rect 7672 13028 7696 13030
rect 7752 13028 7776 13030
rect 7832 13028 7856 13030
rect 7912 13028 7918 13030
rect 7610 13019 7918 13028
rect 7484 12940 7604 12968
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 6950 12540 7258 12549
rect 6950 12538 6956 12540
rect 7012 12538 7036 12540
rect 7092 12538 7116 12540
rect 7172 12538 7196 12540
rect 7252 12538 7258 12540
rect 7012 12486 7014 12538
rect 7194 12486 7196 12538
rect 6950 12484 6956 12486
rect 7012 12484 7036 12486
rect 7092 12484 7116 12486
rect 7172 12484 7196 12486
rect 7252 12484 7258 12486
rect 6950 12475 7258 12484
rect 7104 12232 7156 12238
rect 7288 12232 7340 12238
rect 7104 12174 7156 12180
rect 7194 12200 7250 12209
rect 7116 11558 7144 12174
rect 7288 12174 7340 12180
rect 7194 12135 7196 12144
rect 7248 12135 7250 12144
rect 7196 12106 7248 12112
rect 7300 11898 7328 12174
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7286 11792 7342 11801
rect 7286 11727 7288 11736
rect 7340 11727 7342 11736
rect 7288 11698 7340 11704
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 6950 11452 7258 11461
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 6950 10364 7258 10373
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6950 10299 7258 10308
rect 7300 10146 7328 11290
rect 7208 10118 7328 10146
rect 7208 9602 7236 10118
rect 7286 9752 7342 9761
rect 7286 9687 7288 9696
rect 7340 9687 7342 9696
rect 7288 9658 7340 9664
rect 6920 9580 6972 9586
rect 7208 9574 7328 9602
rect 6920 9522 6972 9528
rect 6932 9489 6960 9522
rect 6918 9480 6974 9489
rect 6918 9415 6974 9424
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 7300 9058 7328 9574
rect 7208 9030 7328 9058
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8498 7052 8774
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7208 8294 7236 9030
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7300 8514 7328 8842
rect 7392 8634 7420 12582
rect 7484 11218 7512 12786
rect 7576 12102 7604 12940
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7748 12640 7800 12646
rect 7746 12608 7748 12617
rect 7800 12608 7802 12617
rect 7746 12543 7802 12552
rect 7746 12336 7802 12345
rect 7746 12271 7802 12280
rect 7656 12232 7708 12238
rect 7760 12220 7788 12271
rect 7708 12192 7788 12220
rect 7656 12174 7708 12180
rect 7852 12170 7880 12786
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7944 12050 7972 12650
rect 8036 12238 8064 13942
rect 8128 13734 8156 14350
rect 8220 14074 8248 14962
rect 8312 14550 8340 15438
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8404 13802 8432 16526
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8392 13796 8444 13802
rect 8392 13738 8444 13744
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8128 12442 8156 13466
rect 8220 12850 8248 13738
rect 8298 13424 8354 13433
rect 8298 13359 8354 13368
rect 8312 12850 8340 13359
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8404 12730 8432 13126
rect 8312 12714 8432 12730
rect 8312 12708 8444 12714
rect 8312 12702 8392 12708
rect 8208 12640 8260 12646
rect 8312 12628 8340 12702
rect 8392 12650 8444 12656
rect 8260 12600 8340 12628
rect 8390 12608 8446 12617
rect 8208 12582 8260 12588
rect 8390 12543 8446 12552
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8300 12368 8352 12374
rect 8404 12345 8432 12543
rect 8300 12310 8352 12316
rect 8390 12336 8446 12345
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8208 12232 8260 12238
rect 8312 12209 8340 12310
rect 8390 12271 8446 12280
rect 8208 12174 8260 12180
rect 8298 12200 8354 12209
rect 8220 12102 8248 12174
rect 8298 12135 8354 12144
rect 8208 12096 8260 12102
rect 7944 12022 8156 12050
rect 8208 12038 8260 12044
rect 7610 11996 7918 12005
rect 7610 11994 7616 11996
rect 7672 11994 7696 11996
rect 7752 11994 7776 11996
rect 7832 11994 7856 11996
rect 7912 11994 7918 11996
rect 7672 11942 7674 11994
rect 7854 11942 7856 11994
rect 7610 11940 7616 11942
rect 7672 11940 7696 11942
rect 7752 11940 7776 11942
rect 7832 11940 7856 11942
rect 7912 11940 7918 11942
rect 7610 11931 7918 11940
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7564 11688 7616 11694
rect 7748 11688 7800 11694
rect 7616 11636 7748 11642
rect 7852 11665 7880 11766
rect 7564 11630 7800 11636
rect 7838 11656 7894 11665
rect 7576 11614 7788 11630
rect 7838 11591 7894 11600
rect 8022 11656 8078 11665
rect 8022 11591 8078 11600
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7576 11098 7604 11494
rect 7668 11286 7696 11494
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7484 11070 7604 11098
rect 7380 8628 7432 8634
rect 7484 8616 7512 11070
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 7562 10296 7618 10305
rect 7562 10231 7618 10240
rect 7576 10130 7604 10231
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 7932 8628 7984 8634
rect 7484 8588 7788 8616
rect 7380 8570 7432 8576
rect 7300 8486 7512 8514
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7116 7478 7144 7890
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7208 7206 7236 8026
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6932 6100 6960 6938
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7024 6322 7052 6870
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6840 6072 6960 6100
rect 6840 5896 6868 6072
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 6840 5868 6960 5896
rect 6734 5808 6790 5817
rect 6734 5743 6790 5752
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6840 4690 6868 5170
rect 6932 5098 6960 5868
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 7300 3738 7328 8366
rect 7484 8294 7512 8486
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7668 8401 7696 8434
rect 7654 8392 7710 8401
rect 7564 8356 7616 8362
rect 7654 8327 7710 8336
rect 7564 8298 7616 8304
rect 7472 8288 7524 8294
rect 7378 8256 7434 8265
rect 7472 8230 7524 8236
rect 7378 8191 7434 8200
rect 7392 5370 7420 8191
rect 7576 7750 7604 8298
rect 7668 8090 7696 8327
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7760 7886 7788 8588
rect 7932 8570 7984 8576
rect 7748 7880 7800 7886
rect 7944 7857 7972 8570
rect 7748 7822 7800 7828
rect 7930 7848 7986 7857
rect 7930 7783 7986 7792
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 7392 2922 7420 5170
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 7484 2446 7512 7142
rect 7852 7002 7880 7346
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 8036 5370 8064 11591
rect 8128 8129 8156 12022
rect 8220 11626 8248 12038
rect 8496 11694 8524 15506
rect 8588 15094 8616 16646
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8588 12186 8616 14486
rect 8680 14006 8708 14826
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8668 13864 8720 13870
rect 8666 13832 8668 13841
rect 8720 13832 8722 13841
rect 8666 13767 8722 13776
rect 8772 13190 8800 16526
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8666 12880 8722 12889
rect 8864 12850 8892 17138
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9048 15609 9076 16390
rect 9034 15600 9090 15609
rect 9034 15535 9090 15544
rect 9140 15473 9168 16526
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 9126 15464 9182 15473
rect 9126 15399 9182 15408
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8956 14822 8984 15098
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 9048 13938 9076 15302
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9140 13841 9168 13874
rect 9126 13832 9182 13841
rect 9126 13767 9182 13776
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 8666 12815 8722 12824
rect 8852 12844 8904 12850
rect 8680 12646 8708 12815
rect 8852 12786 8904 12792
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8850 12744 8906 12753
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8772 12306 8800 12718
rect 8850 12679 8906 12688
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8588 12158 8800 12186
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8298 9888 8354 9897
rect 8114 8120 8170 8129
rect 8114 8055 8170 8064
rect 8220 7970 8248 9862
rect 8298 9823 8354 9832
rect 8312 9722 8340 9823
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8128 7942 8248 7970
rect 8128 5846 8156 7942
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8128 5250 8156 5782
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 8036 5222 8156 5250
rect 7760 5098 7788 5170
rect 8036 5166 8064 5222
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7760 4554 7788 5034
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 8220 2854 8248 7822
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7410 8340 7686
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8404 6866 8432 8842
rect 8496 8634 8524 11630
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8496 7546 8524 7890
rect 8588 7886 8616 8910
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8680 6769 8708 12038
rect 8772 10674 8800 12158
rect 8864 11558 8892 12679
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8666 6760 8722 6769
rect 8666 6695 8722 6704
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8312 5030 8340 5170
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8772 4146 8800 10610
rect 8864 8242 8892 11290
rect 8956 11200 8984 13398
rect 9048 13326 9076 13670
rect 9232 13326 9260 15914
rect 9324 14074 9352 17478
rect 12610 17436 12918 17445
rect 12610 17434 12616 17436
rect 12672 17434 12696 17436
rect 12752 17434 12776 17436
rect 12832 17434 12856 17436
rect 12912 17434 12918 17436
rect 12672 17382 12674 17434
rect 12854 17382 12856 17434
rect 12610 17380 12616 17382
rect 12672 17380 12696 17382
rect 12752 17380 12776 17382
rect 12832 17380 12856 17382
rect 12912 17380 12918 17382
rect 12610 17371 12918 17380
rect 13280 17338 13308 17546
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 13636 17264 13688 17270
rect 13636 17206 13688 17212
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9402 16280 9458 16289
rect 9508 16250 9536 16730
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9402 16215 9458 16224
rect 9496 16244 9548 16250
rect 9416 16182 9444 16215
rect 9496 16186 9548 16192
rect 9404 16176 9456 16182
rect 9404 16118 9456 16124
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9416 15337 9444 15982
rect 9402 15328 9458 15337
rect 9402 15263 9458 15272
rect 9404 15088 9456 15094
rect 9404 15030 9456 15036
rect 9416 14958 9444 15030
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9416 13954 9444 14010
rect 9324 13926 9444 13954
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9324 13308 9352 13926
rect 9404 13320 9456 13326
rect 9324 13280 9404 13308
rect 9232 12458 9260 13262
rect 9048 12430 9260 12458
rect 9048 11354 9076 12430
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 8956 11172 9168 11200
rect 9140 10810 9168 11172
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9048 9518 9076 10746
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8956 8809 8984 8910
rect 8942 8800 8998 8809
rect 8942 8735 8998 8744
rect 8956 8362 8984 8735
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8864 8214 8984 8242
rect 8956 6730 8984 8214
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8864 4622 8892 6258
rect 8956 5137 8984 6666
rect 8942 5128 8998 5137
rect 8942 5063 8998 5072
rect 8956 4690 8984 5063
rect 9048 5030 9076 9454
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 9036 4548 9088 4554
rect 9036 4490 9088 4496
rect 8944 4480 8996 4486
rect 9048 4457 9076 4490
rect 8944 4422 8996 4428
rect 9034 4448 9090 4457
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8850 3632 8906 3641
rect 8850 3567 8906 3576
rect 8864 3058 8892 3567
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8956 2446 8984 4422
rect 9034 4383 9090 4392
rect 9140 3040 9168 10746
rect 9232 7818 9260 11290
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9232 4690 9260 7754
rect 9324 7002 9352 13280
rect 9404 13262 9456 13268
rect 9508 12481 9536 14758
rect 9600 14498 9628 16526
rect 9692 16046 9720 16662
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9784 15473 9812 16934
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9876 16182 9904 16730
rect 10060 16590 10088 17070
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9968 16114 9996 16458
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9770 15464 9826 15473
rect 9770 15399 9826 15408
rect 9678 15192 9734 15201
rect 9678 15127 9680 15136
rect 9732 15127 9734 15136
rect 9680 15098 9732 15104
rect 9784 15042 9812 15399
rect 9692 15026 9812 15042
rect 9680 15020 9812 15026
rect 9732 15014 9812 15020
rect 9680 14962 9732 14968
rect 9772 14952 9824 14958
rect 9770 14920 9772 14929
rect 9824 14920 9826 14929
rect 9680 14884 9732 14890
rect 9770 14855 9826 14864
rect 9680 14826 9732 14832
rect 9692 14793 9720 14826
rect 9678 14784 9734 14793
rect 9678 14719 9734 14728
rect 9678 14648 9734 14657
rect 9678 14583 9680 14592
rect 9732 14583 9734 14592
rect 9680 14554 9732 14560
rect 9784 14521 9812 14855
rect 9770 14512 9826 14521
rect 9600 14470 9720 14498
rect 9586 14376 9642 14385
rect 9586 14311 9642 14320
rect 9600 14278 9628 14311
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9692 14090 9720 14470
rect 9770 14447 9826 14456
rect 9600 14074 9720 14090
rect 9588 14068 9720 14074
rect 9640 14062 9720 14068
rect 9588 14010 9640 14016
rect 9772 13320 9824 13326
rect 9586 13288 9642 13297
rect 9772 13262 9824 13268
rect 9586 13223 9588 13232
rect 9640 13223 9642 13232
rect 9588 13194 9640 13200
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9494 12472 9550 12481
rect 9494 12407 9550 12416
rect 9404 12232 9456 12238
rect 9600 12220 9628 12786
rect 9678 12744 9734 12753
rect 9678 12679 9734 12688
rect 9692 12442 9720 12679
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9678 12336 9734 12345
rect 9678 12271 9680 12280
rect 9732 12271 9734 12280
rect 9680 12242 9732 12248
rect 9456 12192 9628 12220
rect 9404 12174 9456 12180
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9324 5642 9352 6938
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4690 9352 4966
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4282 9352 4422
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9324 3534 9352 4218
rect 9416 3942 9444 12174
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9508 11801 9536 12038
rect 9588 11824 9640 11830
rect 9494 11792 9550 11801
rect 9588 11766 9640 11772
rect 9494 11727 9550 11736
rect 9600 10996 9628 11766
rect 9508 10968 9628 10996
rect 9508 6322 9536 10968
rect 9586 9616 9642 9625
rect 9692 9586 9720 12038
rect 9784 10169 9812 13262
rect 9876 12889 9904 15846
rect 9862 12880 9918 12889
rect 9862 12815 9918 12824
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9876 11150 9904 12106
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9770 10160 9826 10169
rect 9770 10095 9826 10104
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9586 9551 9642 9560
rect 9680 9580 9732 9586
rect 9600 8566 9628 9551
rect 9680 9522 9732 9528
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9784 8401 9812 9930
rect 9770 8392 9826 8401
rect 9680 8356 9732 8362
rect 9770 8327 9826 8336
rect 9680 8298 9732 8304
rect 9692 6458 9720 8298
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9784 6798 9812 8230
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 6458 9812 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9876 4282 9904 11086
rect 9968 10606 9996 16050
rect 10060 15745 10088 16050
rect 10046 15736 10102 15745
rect 10046 15671 10102 15680
rect 10152 15586 10180 16390
rect 10060 15558 10180 15586
rect 10060 13938 10088 15558
rect 10138 15056 10194 15065
rect 10138 14991 10194 15000
rect 10152 14958 10180 14991
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10244 14770 10272 17002
rect 10324 16584 10376 16590
rect 10322 16552 10324 16561
rect 10376 16552 10378 16561
rect 10322 16487 10378 16496
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 15201 10364 16390
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 15337 10456 15438
rect 10414 15328 10470 15337
rect 10414 15263 10470 15272
rect 10322 15192 10378 15201
rect 10322 15127 10378 15136
rect 10520 14890 10548 17206
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10600 16516 10652 16522
rect 10600 16458 10652 16464
rect 10612 15337 10640 16458
rect 10704 15570 10732 16594
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10690 15464 10746 15473
rect 10690 15399 10746 15408
rect 10598 15328 10654 15337
rect 10598 15263 10654 15272
rect 10704 15162 10732 15399
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10612 14793 10640 14962
rect 10598 14784 10654 14793
rect 10244 14742 10456 14770
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10152 13977 10180 14554
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10244 14074 10272 14418
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10138 13968 10194 13977
rect 10048 13932 10100 13938
rect 10138 13903 10194 13912
rect 10048 13874 10100 13880
rect 10060 13530 10088 13874
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 9722 9996 10542
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 10060 9654 10088 13466
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10060 8498 10088 9590
rect 10048 8492 10100 8498
rect 9968 8452 10048 8480
rect 9968 6798 9996 8452
rect 10048 8434 10100 8440
rect 10152 7954 10180 12378
rect 10244 11694 10272 14010
rect 10322 13968 10378 13977
rect 10322 13903 10378 13912
rect 10336 12986 10364 13903
rect 10428 12986 10456 14742
rect 10598 14719 10654 14728
rect 10506 14648 10562 14657
rect 10506 14583 10562 14592
rect 10520 14482 10548 14583
rect 10598 14512 10654 14521
rect 10508 14476 10560 14482
rect 10598 14447 10654 14456
rect 10508 14418 10560 14424
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10336 12322 10364 12786
rect 10428 12442 10456 12922
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10336 12294 10456 12322
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10336 9761 10364 12174
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 6186 9996 6598
rect 10060 6254 10088 6734
rect 10152 6390 10180 6802
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9954 4312 10010 4321
rect 9864 4276 9916 4282
rect 10152 4282 10180 6326
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 4690 10272 6054
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 9954 4247 10010 4256
rect 10140 4276 10192 4282
rect 9864 4218 9916 4224
rect 9968 4214 9996 4247
rect 10140 4218 10192 4224
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10152 4049 10180 4082
rect 10138 4040 10194 4049
rect 10336 4010 10364 9687
rect 10428 9450 10456 12294
rect 10520 12102 10548 12786
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10506 11928 10562 11937
rect 10506 11863 10562 11872
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10520 8362 10548 11863
rect 10612 11762 10640 14447
rect 10704 12850 10732 15098
rect 10796 13462 10824 16934
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10796 12434 10824 13398
rect 10704 12406 10824 12434
rect 10704 12170 10732 12406
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10138 3975 10194 3984
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9600 3194 9628 3470
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 10520 3058 10548 8298
rect 10612 6458 10640 9998
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10704 6390 10732 12106
rect 10888 11082 10916 16526
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10980 15706 11008 15982
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10980 15337 11008 15506
rect 10966 15328 11022 15337
rect 10966 15263 11022 15272
rect 10966 15192 11022 15201
rect 10966 15127 11022 15136
rect 10980 14278 11008 15127
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10980 13190 11008 13330
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 11072 12730 11100 15846
rect 10980 12702 11100 12730
rect 10980 11914 11008 12702
rect 11058 12608 11114 12617
rect 11058 12543 11114 12552
rect 11072 12102 11100 12543
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10980 11886 11100 11914
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10980 10996 11008 11494
rect 11072 11150 11100 11886
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10980 10968 11100 10996
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10704 6118 10732 6326
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 9220 3052 9272 3058
rect 9140 3012 9220 3040
rect 9220 2994 9272 3000
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 9126 2680 9182 2689
rect 9126 2615 9182 2624
rect 9140 2446 9168 2615
rect 10704 2514 10732 2994
rect 10796 2582 10824 9522
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10888 7002 10916 8434
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10888 5302 10916 5646
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10980 3398 11008 9862
rect 11072 6798 11100 10968
rect 11164 10198 11192 16390
rect 11256 12617 11284 16730
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11242 12608 11298 12617
rect 11242 12543 11298 12552
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11164 7478 11192 8570
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11164 6730 11192 7278
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11072 5098 11100 5306
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 11072 4622 11100 5034
rect 11164 5030 11192 6666
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11150 4856 11206 4865
rect 11150 4791 11206 4800
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11164 4554 11192 4791
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10966 3224 11022 3233
rect 10966 3159 10968 3168
rect 11020 3159 11022 3168
rect 10968 3130 11020 3136
rect 11072 2650 11100 4150
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11164 3058 11192 3538
rect 11256 3466 11284 12378
rect 11348 9994 11376 15982
rect 11428 15972 11480 15978
rect 11428 15914 11480 15920
rect 11440 15706 11468 15914
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11426 15464 11482 15473
rect 11426 15399 11482 15408
rect 11440 14249 11468 15399
rect 11426 14240 11482 14249
rect 11426 14175 11482 14184
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11440 13394 11468 13806
rect 11532 13734 11560 16186
rect 11808 15910 11836 17002
rect 11950 16892 12258 16901
rect 11950 16890 11956 16892
rect 12012 16890 12036 16892
rect 12092 16890 12116 16892
rect 12172 16890 12196 16892
rect 12252 16890 12258 16892
rect 12012 16838 12014 16890
rect 12194 16838 12196 16890
rect 11950 16836 11956 16838
rect 12012 16836 12036 16838
rect 12092 16836 12116 16838
rect 12172 16836 12196 16838
rect 12252 16836 12258 16838
rect 11950 16827 12258 16836
rect 13648 16658 13676 17206
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 11978 16280 12034 16289
rect 11978 16215 12034 16224
rect 11992 16182 12020 16215
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 12254 16144 12310 16153
rect 12310 16102 12388 16130
rect 12254 16079 12310 16088
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11950 15804 12258 15813
rect 11950 15802 11956 15804
rect 12012 15802 12036 15804
rect 12092 15802 12116 15804
rect 12172 15802 12196 15804
rect 12252 15802 12258 15804
rect 12012 15750 12014 15802
rect 12194 15750 12196 15802
rect 11950 15748 11956 15750
rect 12012 15748 12036 15750
rect 12092 15748 12116 15750
rect 12172 15748 12196 15750
rect 12252 15748 12258 15750
rect 11950 15739 12258 15748
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11440 12306 11468 12650
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11624 12238 11652 14962
rect 12360 14793 12388 16102
rect 12346 14784 12402 14793
rect 11950 14716 12258 14725
rect 12346 14719 12402 14728
rect 11950 14714 11956 14716
rect 12012 14714 12036 14716
rect 12092 14714 12116 14716
rect 12172 14714 12196 14716
rect 12252 14714 12258 14716
rect 12012 14662 12014 14714
rect 12194 14662 12196 14714
rect 11950 14660 11956 14662
rect 12012 14660 12036 14662
rect 12092 14660 12116 14662
rect 12172 14660 12196 14662
rect 12252 14660 12258 14662
rect 11950 14651 12258 14660
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11716 12442 11744 14282
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 11950 13628 12258 13637
rect 11950 13626 11956 13628
rect 12012 13626 12036 13628
rect 12092 13626 12116 13628
rect 12172 13626 12196 13628
rect 12252 13626 12258 13628
rect 12012 13574 12014 13626
rect 12194 13574 12196 13626
rect 11950 13572 11956 13574
rect 12012 13572 12036 13574
rect 12092 13572 12116 13574
rect 12172 13572 12196 13574
rect 12252 13572 12258 13574
rect 11950 13563 12258 13572
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12268 12850 12296 13330
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11702 12336 11758 12345
rect 11702 12271 11758 12280
rect 11716 12238 11744 12271
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11428 12096 11480 12102
rect 11624 12084 11652 12174
rect 11624 12056 11744 12084
rect 11428 12038 11480 12044
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 11440 9874 11468 12038
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11532 11393 11560 11494
rect 11518 11384 11574 11393
rect 11518 11319 11574 11328
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11348 9846 11468 9874
rect 11348 8634 11376 9846
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11532 8498 11560 11086
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 3534 11376 7142
rect 11440 5778 11468 7414
rect 11532 6730 11560 8026
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11440 3058 11468 4966
rect 11624 4622 11652 11562
rect 11716 9489 11744 12056
rect 11808 11150 11836 12786
rect 11950 12540 12258 12549
rect 11950 12538 11956 12540
rect 12012 12538 12036 12540
rect 12092 12538 12116 12540
rect 12172 12538 12196 12540
rect 12252 12538 12258 12540
rect 12012 12486 12014 12538
rect 12194 12486 12196 12538
rect 11950 12484 11956 12486
rect 12012 12484 12036 12486
rect 12092 12484 12116 12486
rect 12172 12484 12196 12486
rect 12252 12484 12258 12486
rect 11950 12475 12258 12484
rect 11888 12436 11940 12442
rect 12360 12434 12388 13942
rect 11888 12378 11940 12384
rect 12084 12406 12388 12434
rect 11900 12306 11928 12378
rect 11978 12336 12034 12345
rect 11888 12300 11940 12306
rect 11978 12271 12034 12280
rect 11888 12242 11940 12248
rect 11886 11928 11942 11937
rect 11886 11863 11942 11872
rect 11900 11762 11928 11863
rect 11992 11830 12020 12271
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 12084 11558 12112 12406
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12176 11626 12204 12174
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11950 11452 12258 11461
rect 11950 11450 11956 11452
rect 12012 11450 12036 11452
rect 12092 11450 12116 11452
rect 12172 11450 12196 11452
rect 12252 11450 12258 11452
rect 12012 11398 12014 11450
rect 12194 11398 12196 11450
rect 11950 11396 11956 11398
rect 12012 11396 12036 11398
rect 12092 11396 12116 11398
rect 12172 11396 12196 11398
rect 12252 11396 12258 11398
rect 11950 11387 12258 11396
rect 12360 11150 12388 12242
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 11794 10840 11850 10849
rect 11794 10775 11850 10784
rect 11808 10470 11836 10775
rect 12268 10674 12296 11086
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11702 9480 11758 9489
rect 11702 9415 11758 9424
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11716 8809 11744 8978
rect 11702 8800 11758 8809
rect 11702 8735 11758 8744
rect 11716 5098 11744 8735
rect 11808 6254 11836 10406
rect 11950 10364 12258 10373
rect 11950 10362 11956 10364
rect 12012 10362 12036 10364
rect 12092 10362 12116 10364
rect 12172 10362 12196 10364
rect 12252 10362 12258 10364
rect 12012 10310 12014 10362
rect 12194 10310 12196 10362
rect 11950 10308 11956 10310
rect 12012 10308 12036 10310
rect 12092 10308 12116 10310
rect 12172 10308 12196 10310
rect 12252 10308 12258 10310
rect 11950 10299 12258 10308
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11900 9722 11928 9998
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11950 9276 12258 9285
rect 11950 9274 11956 9276
rect 12012 9274 12036 9276
rect 12092 9274 12116 9276
rect 12172 9274 12196 9276
rect 12252 9274 12258 9276
rect 12012 9222 12014 9274
rect 12194 9222 12196 9274
rect 11950 9220 11956 9222
rect 12012 9220 12036 9222
rect 12092 9220 12116 9222
rect 12172 9220 12196 9222
rect 12252 9220 12258 9222
rect 11950 9211 12258 9220
rect 12360 9042 12388 11086
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12452 8634 12480 16458
rect 13280 16425 13308 16458
rect 13266 16416 13322 16425
rect 12610 16348 12918 16357
rect 13266 16351 13322 16360
rect 12610 16346 12616 16348
rect 12672 16346 12696 16348
rect 12752 16346 12776 16348
rect 12832 16346 12856 16348
rect 12912 16346 12918 16348
rect 12672 16294 12674 16346
rect 12854 16294 12856 16346
rect 12610 16292 12616 16294
rect 12672 16292 12696 16294
rect 12752 16292 12776 16294
rect 12832 16292 12856 16294
rect 12912 16292 12918 16294
rect 12610 16283 12918 16292
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 12992 16108 13044 16114
rect 13188 16096 13216 16186
rect 13268 16108 13320 16114
rect 13188 16068 13268 16096
rect 12992 16050 13044 16056
rect 13268 16050 13320 16056
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12912 15434 12940 15982
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12530 14648 12586 14657
rect 12636 14618 12664 15030
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12530 14583 12586 14592
rect 12624 14612 12676 14618
rect 12544 14006 12572 14583
rect 12624 14554 12676 14560
rect 12912 14550 12940 14894
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12532 13728 12584 13734
rect 13004 13705 13032 16050
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 12532 13670 12584 13676
rect 12990 13696 13046 13705
rect 12544 13326 12572 13670
rect 12990 13631 13046 13640
rect 13096 13546 13124 14486
rect 13004 13518 13124 13546
rect 13188 13530 13216 15438
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 13176 13524 13228 13530
rect 12714 13424 12770 13433
rect 12714 13359 12770 13368
rect 12728 13326 12756 13359
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 13004 12714 13032 13518
rect 13176 13466 13228 13472
rect 13280 13410 13308 15370
rect 13464 14550 13492 16050
rect 13634 16008 13690 16017
rect 13634 15943 13690 15952
rect 13542 15600 13598 15609
rect 13542 15535 13544 15544
rect 13596 15535 13598 15544
rect 13544 15506 13596 15512
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14618 13584 14758
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13372 14006 13400 14418
rect 13360 14000 13412 14006
rect 13648 13954 13676 15943
rect 13740 15722 13768 17206
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 14464 17128 14516 17134
rect 14094 17096 14150 17105
rect 14464 17070 14516 17076
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 14094 17031 14150 17040
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13740 15694 13860 15722
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13740 15094 13768 15506
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13832 14362 13860 15694
rect 13360 13942 13412 13948
rect 13556 13926 13676 13954
rect 13740 14334 13860 14362
rect 13556 13734 13584 13926
rect 13636 13864 13688 13870
rect 13634 13832 13636 13841
rect 13688 13832 13690 13841
rect 13634 13767 13690 13776
rect 13544 13728 13596 13734
rect 13450 13696 13506 13705
rect 13544 13670 13596 13676
rect 13450 13631 13506 13640
rect 13188 13382 13308 13410
rect 13360 13388 13412 13394
rect 13082 13016 13138 13025
rect 13082 12951 13084 12960
rect 13136 12951 13138 12960
rect 13084 12922 13136 12928
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12544 11218 12572 12582
rect 12622 12472 12678 12481
rect 12622 12407 12678 12416
rect 12636 12238 12664 12407
rect 12992 12368 13044 12374
rect 12990 12336 12992 12345
rect 13044 12336 13046 12345
rect 12990 12271 13046 12280
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12624 11552 12676 11558
rect 12728 11529 12756 11834
rect 13004 11665 13032 12174
rect 13188 11914 13216 13382
rect 13360 13330 13412 13336
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13280 12345 13308 12922
rect 13266 12336 13322 12345
rect 13266 12271 13322 12280
rect 13096 11898 13216 11914
rect 13084 11892 13216 11898
rect 13136 11886 13216 11892
rect 13084 11834 13136 11840
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 12990 11656 13046 11665
rect 12990 11591 13046 11600
rect 12992 11552 13044 11558
rect 12624 11494 12676 11500
rect 12714 11520 12770 11529
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12636 11014 12664 11494
rect 12992 11494 13044 11500
rect 12714 11455 12770 11464
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12610 10843 12918 10852
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12544 8498 12572 10610
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12636 10130 12664 10474
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 8294 12572 8434
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 11950 8188 12258 8197
rect 11950 8186 11956 8188
rect 12012 8186 12036 8188
rect 12092 8186 12116 8188
rect 12172 8186 12196 8188
rect 12252 8186 12258 8188
rect 12012 8134 12014 8186
rect 12194 8134 12196 8186
rect 11950 8132 11956 8134
rect 12012 8132 12036 8134
rect 12092 8132 12116 8134
rect 12172 8132 12196 8134
rect 12252 8132 12258 8134
rect 11950 8123 12258 8132
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 11950 7100 12258 7109
rect 11950 7098 11956 7100
rect 12012 7098 12036 7100
rect 12092 7098 12116 7100
rect 12172 7098 12196 7100
rect 12252 7098 12258 7100
rect 12012 7046 12014 7098
rect 12194 7046 12196 7098
rect 11950 7044 11956 7046
rect 12012 7044 12036 7046
rect 12092 7044 12116 7046
rect 12172 7044 12196 7046
rect 12252 7044 12258 7046
rect 11950 7035 12258 7044
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12360 6730 12388 6802
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12452 6610 12480 7414
rect 12530 6896 12586 6905
rect 12530 6831 12586 6840
rect 12544 6798 12572 6831
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12452 6582 12572 6610
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 11950 6012 12258 6021
rect 11950 6010 11956 6012
rect 12012 6010 12036 6012
rect 12092 6010 12116 6012
rect 12172 6010 12196 6012
rect 12252 6010 12258 6012
rect 12012 5958 12014 6010
rect 12194 5958 12196 6010
rect 11950 5956 11956 5958
rect 12012 5956 12036 5958
rect 12092 5956 12116 5958
rect 12172 5956 12196 5958
rect 12252 5956 12258 5958
rect 11950 5947 12258 5956
rect 12360 5710 12388 6190
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12254 5264 12310 5273
rect 12254 5199 12256 5208
rect 12308 5199 12310 5208
rect 12256 5170 12308 5176
rect 11704 5092 11756 5098
rect 11704 5034 11756 5040
rect 11950 4924 12258 4933
rect 11950 4922 11956 4924
rect 12012 4922 12036 4924
rect 12092 4922 12116 4924
rect 12172 4922 12196 4924
rect 12252 4922 12258 4924
rect 12012 4870 12014 4922
rect 12194 4870 12196 4922
rect 11950 4868 11956 4870
rect 12012 4868 12036 4870
rect 12092 4868 12116 4870
rect 12172 4868 12196 4870
rect 12252 4868 12258 4870
rect 11950 4859 12258 4868
rect 12452 4758 12480 6054
rect 12072 4752 12124 4758
rect 12070 4720 12072 4729
rect 12440 4752 12492 4758
rect 12124 4720 12126 4729
rect 12070 4655 12126 4664
rect 12254 4720 12310 4729
rect 12440 4694 12492 4700
rect 12544 4690 12572 6582
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 13004 5302 13032 11494
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13096 5556 13124 9114
rect 13188 5914 13216 11766
rect 13280 11558 13308 12271
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13280 10606 13308 10950
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13280 9178 13308 10542
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13266 8936 13322 8945
rect 13266 8871 13322 8880
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13176 5568 13228 5574
rect 13096 5528 13176 5556
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 13096 4758 13124 5528
rect 13176 5510 13228 5516
rect 13280 5234 13308 8871
rect 13372 6186 13400 13330
rect 13464 12481 13492 13631
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13556 12866 13584 13466
rect 13740 13410 13768 14334
rect 13820 13864 13872 13870
rect 13818 13832 13820 13841
rect 13872 13832 13874 13841
rect 13818 13767 13874 13776
rect 13648 13382 13768 13410
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13648 12986 13676 13382
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13556 12838 13676 12866
rect 13450 12472 13506 12481
rect 13450 12407 13506 12416
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13452 12096 13504 12102
rect 13450 12064 13452 12073
rect 13504 12064 13506 12073
rect 13450 11999 13506 12008
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 13464 5234 13492 11999
rect 13556 5710 13584 12174
rect 13648 11830 13676 12838
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13648 10130 13676 10610
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13740 9722 13768 13262
rect 13832 12850 13860 13398
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13924 12306 13952 16662
rect 14108 15706 14136 17031
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14186 16552 14242 16561
rect 14186 16487 14188 16496
rect 14240 16487 14242 16496
rect 14188 16458 14240 16464
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14108 14958 14136 15438
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14096 14952 14148 14958
rect 14016 14912 14096 14940
rect 14016 13870 14044 14912
rect 14096 14894 14148 14900
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14108 13394 14136 14486
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14002 12880 14058 12889
rect 14002 12815 14058 12824
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13818 10704 13874 10713
rect 13818 10639 13820 10648
rect 13872 10639 13874 10648
rect 13820 10610 13872 10616
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13740 8430 13768 9658
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13648 7478 13676 7686
rect 13636 7472 13688 7478
rect 13636 7414 13688 7420
rect 13832 7410 13860 9930
rect 13924 7546 13952 12038
rect 14016 10470 14044 12815
rect 14108 12306 14136 13126
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14108 11132 14136 11834
rect 14200 11762 14228 14962
rect 14292 14657 14320 16594
rect 14476 16590 14504 17070
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14660 16658 14688 16934
rect 15212 16697 15240 17070
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15672 16794 15700 17002
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15198 16688 15254 16697
rect 14648 16652 14700 16658
rect 15198 16623 15254 16632
rect 14648 16594 14700 16600
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 14372 14952 14424 14958
rect 14370 14920 14372 14929
rect 14424 14920 14426 14929
rect 14370 14855 14426 14864
rect 14476 14822 14504 16526
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14568 15026 14596 16050
rect 14936 16046 14964 16390
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14278 14648 14334 14657
rect 14278 14583 14334 14592
rect 14292 12986 14320 14583
rect 14554 14512 14610 14521
rect 14554 14447 14610 14456
rect 14568 13938 14596 14447
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14384 12918 14412 13874
rect 14556 13320 14608 13326
rect 14554 13288 14556 13297
rect 14608 13288 14610 13297
rect 14464 13252 14516 13258
rect 14554 13223 14610 13232
rect 14464 13194 14516 13200
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14292 12238 14320 12650
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14292 11830 14320 12174
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14200 11393 14228 11698
rect 14384 11558 14412 12242
rect 14476 12238 14504 13194
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14186 11384 14242 11393
rect 14186 11319 14242 11328
rect 14188 11144 14240 11150
rect 14108 11104 14188 11132
rect 14108 11014 14136 11104
rect 14188 11086 14240 11092
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14188 10668 14240 10674
rect 14240 10628 14320 10656
rect 14188 10610 14240 10616
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13818 6896 13874 6905
rect 13818 6831 13874 6840
rect 13726 6488 13782 6497
rect 13726 6423 13782 6432
rect 13740 6390 13768 6423
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13832 6254 13860 6831
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13818 5944 13874 5953
rect 13818 5879 13874 5888
rect 13832 5846 13860 5879
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13556 5574 13584 5646
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13176 5160 13228 5166
rect 13174 5128 13176 5137
rect 13228 5128 13230 5137
rect 13174 5063 13230 5072
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12254 4655 12310 4664
rect 12532 4684 12584 4690
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 12268 4185 12296 4655
rect 12532 4626 12584 4632
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12360 4457 12388 4490
rect 12346 4448 12402 4457
rect 12346 4383 12402 4392
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 12254 4176 12310 4185
rect 12254 4111 12310 4120
rect 12346 4040 12402 4049
rect 12346 3975 12348 3984
rect 12400 3975 12402 3984
rect 12348 3946 12400 3952
rect 11950 3836 12258 3845
rect 11950 3834 11956 3836
rect 12012 3834 12036 3836
rect 12092 3834 12116 3836
rect 12172 3834 12196 3836
rect 12252 3834 12258 3836
rect 12012 3782 12014 3834
rect 12194 3782 12196 3834
rect 11950 3780 11956 3782
rect 12012 3780 12036 3782
rect 12092 3780 12116 3782
rect 12172 3780 12196 3782
rect 12252 3780 12258 3782
rect 11950 3771 12258 3780
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12176 3058 12204 3470
rect 12360 3126 12388 3946
rect 13096 3534 13124 4694
rect 13464 3670 13492 5170
rect 13740 4826 13768 5170
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12544 3058 12572 3334
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 11950 2748 12258 2757
rect 11950 2746 11956 2748
rect 12012 2746 12036 2748
rect 12092 2746 12116 2748
rect 12172 2746 12196 2748
rect 12252 2746 12258 2748
rect 12012 2694 12014 2746
rect 12194 2694 12196 2746
rect 11950 2692 11956 2694
rect 12012 2692 12036 2694
rect 12092 2692 12116 2694
rect 12172 2692 12196 2694
rect 12252 2692 12258 2694
rect 11950 2683 12258 2692
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 13740 2378 13768 4762
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13832 4486 13860 4626
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13924 3126 13952 7482
rect 14016 7342 14044 9998
rect 14292 9926 14320 10628
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14094 8392 14150 8401
rect 14200 8378 14228 8978
rect 14292 8514 14320 9862
rect 14384 8634 14412 11494
rect 14476 11014 14504 12174
rect 14568 11830 14596 12922
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14292 8486 14412 8514
rect 14200 8350 14320 8378
rect 14094 8327 14150 8336
rect 14108 7410 14136 8327
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14200 7410 14228 7890
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14016 6866 14044 7278
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14016 4486 14044 6598
rect 14200 5794 14228 7346
rect 14292 6322 14320 8350
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14200 5766 14320 5794
rect 14292 5710 14320 5766
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14094 5264 14150 5273
rect 14094 5199 14150 5208
rect 14108 4826 14136 5199
rect 14384 4978 14412 8486
rect 14476 8430 14504 10950
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14464 8288 14516 8294
rect 14568 8242 14596 11222
rect 14660 11082 14688 15846
rect 14936 15502 14964 15982
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14830 15056 14886 15065
rect 14830 14991 14886 15000
rect 14844 14890 14872 14991
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14660 8838 14688 10542
rect 14752 8974 14780 14758
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14936 14278 14964 14554
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14844 13705 14872 13874
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 15028 13818 15056 16526
rect 14830 13696 14886 13705
rect 14830 13631 14886 13640
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14844 11626 14872 13262
rect 14936 13172 14964 13806
rect 15028 13802 15148 13818
rect 15028 13796 15160 13802
rect 15028 13790 15108 13796
rect 15108 13738 15160 13744
rect 15212 13462 15240 16526
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15396 15434 15424 16458
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15488 15978 15516 16186
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15488 15502 15516 15914
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 14936 13144 15056 13172
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 14830 11248 14886 11257
rect 14830 11183 14832 11192
rect 14884 11183 14886 11192
rect 14832 11154 14884 11160
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14516 8236 14596 8242
rect 14464 8230 14596 8236
rect 14476 8214 14596 8230
rect 14476 7206 14504 8214
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 5114 14504 7142
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14568 5302 14596 5510
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 14476 5086 14596 5114
rect 14384 4950 14504 4978
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14476 4622 14504 4950
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3505 14412 3878
rect 14476 3602 14504 4558
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14370 3496 14426 3505
rect 14370 3431 14426 3440
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 14568 3058 14596 5086
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14660 2990 14688 8774
rect 14844 8498 14872 11018
rect 14936 10606 14964 12786
rect 15028 11626 15056 13144
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15108 11824 15160 11830
rect 15108 11766 15160 11772
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 15028 11218 15056 11562
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15120 10985 15148 11766
rect 15106 10976 15162 10985
rect 15106 10911 15162 10920
rect 15212 10826 15240 12310
rect 15304 11354 15332 13874
rect 15396 11898 15424 15370
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 12442 15516 13670
rect 15580 13326 15608 13738
rect 15672 13569 15700 14214
rect 15658 13560 15714 13569
rect 15658 13495 15714 13504
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15396 11121 15424 11698
rect 15382 11112 15438 11121
rect 15382 11047 15438 11056
rect 15108 10804 15160 10810
rect 15212 10798 15332 10826
rect 15108 10746 15160 10752
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15028 10305 15056 10610
rect 15014 10296 15070 10305
rect 15014 10231 15070 10240
rect 14924 10192 14976 10198
rect 14924 10134 14976 10140
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14752 4214 14780 8366
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14844 5914 14872 7686
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14830 5808 14886 5817
rect 14830 5743 14886 5752
rect 14844 5710 14872 5743
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14936 4486 14964 10134
rect 15120 10062 15148 10746
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15212 10062 15240 10678
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15198 9752 15254 9761
rect 15198 9687 15254 9696
rect 15212 9586 15240 9687
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15028 8838 15056 9386
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15120 8945 15148 9114
rect 15200 8968 15252 8974
rect 15106 8936 15162 8945
rect 15200 8910 15252 8916
rect 15106 8871 15162 8880
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 15212 8537 15240 8910
rect 15198 8528 15254 8537
rect 15198 8463 15254 8472
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15106 6896 15162 6905
rect 15106 6831 15162 6840
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 15028 3126 15056 5850
rect 15120 4214 15148 6831
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 15120 3738 15148 4150
rect 15212 4146 15240 7142
rect 15304 5234 15332 10798
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15396 10198 15424 10542
rect 15384 10192 15436 10198
rect 15384 10134 15436 10140
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15396 9722 15424 9930
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15396 9042 15424 9522
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15382 8256 15438 8265
rect 15382 8191 15438 8200
rect 15396 5710 15424 8191
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15396 4729 15424 5170
rect 15382 4720 15438 4729
rect 15382 4655 15438 4664
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 15304 2582 15332 4082
rect 15488 3602 15516 12106
rect 15672 11914 15700 13330
rect 15764 12434 15792 14418
rect 15856 13433 15884 15846
rect 15842 13424 15898 13433
rect 15842 13359 15898 13368
rect 15764 12406 15884 12434
rect 15672 11886 15792 11914
rect 15658 11520 15714 11529
rect 15658 11455 15714 11464
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15580 2650 15608 11222
rect 15672 8498 15700 11455
rect 15764 9761 15792 11886
rect 15856 11694 15884 12406
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15750 9752 15806 9761
rect 15750 9687 15806 9696
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15764 9110 15792 9522
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15658 7304 15714 7313
rect 15658 7239 15714 7248
rect 15672 6730 15700 7239
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15856 6186 15884 11630
rect 15948 11218 15976 16390
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15934 11112 15990 11121
rect 15934 11047 15990 11056
rect 15948 9466 15976 11047
rect 16040 9722 16068 13262
rect 16132 13025 16160 14962
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16118 13016 16174 13025
rect 16118 12951 16174 12960
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 11082 16160 11494
rect 16224 11354 16252 13330
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16210 11112 16266 11121
rect 16120 11076 16172 11082
rect 16210 11047 16266 11056
rect 16120 11018 16172 11024
rect 16224 10962 16252 11047
rect 16132 10934 16252 10962
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 15948 9438 16068 9466
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15948 5778 15976 9318
rect 16040 6934 16068 9438
rect 16132 6934 16160 10934
rect 16316 9625 16344 12378
rect 16408 11665 16436 17138
rect 16592 15502 16620 17546
rect 17610 17436 17918 17445
rect 17610 17434 17616 17436
rect 17672 17434 17696 17436
rect 17752 17434 17776 17436
rect 17832 17434 17856 17436
rect 17912 17434 17918 17436
rect 17672 17382 17674 17434
rect 17854 17382 17856 17434
rect 17610 17380 17616 17382
rect 17672 17380 17696 17382
rect 17752 17380 17776 17382
rect 17832 17380 17856 17382
rect 17912 17380 17918 17382
rect 17610 17371 17918 17380
rect 17972 17338 18000 17598
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 16950 16892 17258 16901
rect 16950 16890 16956 16892
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17252 16890 17258 16892
rect 17012 16838 17014 16890
rect 17194 16838 17196 16890
rect 16950 16836 16956 16838
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 17252 16836 17258 16838
rect 16950 16827 17258 16836
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16592 14906 16620 15438
rect 16500 14878 16620 14906
rect 16500 12322 16528 14878
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 12442 16620 14758
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16500 12294 16620 12322
rect 16394 11656 16450 11665
rect 16394 11591 16450 11600
rect 16408 11121 16436 11591
rect 16394 11112 16450 11121
rect 16394 11047 16450 11056
rect 16486 10568 16542 10577
rect 16486 10503 16542 10512
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16302 9616 16358 9625
rect 16302 9551 16358 9560
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 8022 16344 9318
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16316 7002 16344 7278
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16028 6928 16080 6934
rect 16028 6870 16080 6876
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16118 6760 16174 6769
rect 16118 6695 16174 6704
rect 16212 6724 16264 6730
rect 16132 6254 16160 6695
rect 16212 6666 16264 6672
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16224 6186 16252 6666
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16224 5370 16252 5510
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16316 4826 16344 6258
rect 16408 5302 16436 9930
rect 16500 6322 16528 10503
rect 16592 10198 16620 12294
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16578 10024 16634 10033
rect 16578 9959 16634 9968
rect 16592 9722 16620 9959
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16488 6180 16540 6186
rect 16488 6122 16540 6128
rect 16500 5778 16528 6122
rect 16592 5914 16620 9522
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16592 5658 16620 5850
rect 16500 5642 16620 5658
rect 16488 5636 16620 5642
rect 16540 5630 16620 5636
rect 16488 5578 16540 5584
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 16684 4826 16712 16526
rect 16776 15042 16804 16662
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16868 15609 16896 16526
rect 16960 16017 16988 16526
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 16946 16008 17002 16017
rect 16946 15943 17002 15952
rect 16950 15804 17258 15813
rect 16950 15802 16956 15804
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17252 15802 17258 15804
rect 17012 15750 17014 15802
rect 17194 15750 17196 15802
rect 16950 15748 16956 15750
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 17252 15748 17258 15750
rect 16950 15739 17258 15748
rect 16854 15600 16910 15609
rect 16854 15535 16910 15544
rect 17132 15496 17184 15502
rect 16854 15464 16910 15473
rect 17132 15438 17184 15444
rect 16854 15399 16856 15408
rect 16908 15399 16910 15408
rect 16856 15370 16908 15376
rect 17144 15094 17172 15438
rect 17132 15088 17184 15094
rect 16776 15014 16896 15042
rect 17132 15030 17184 15036
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16776 14793 16804 14894
rect 16762 14784 16818 14793
rect 16762 14719 16818 14728
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16776 12889 16804 14282
rect 16762 12880 16818 12889
rect 16762 12815 16818 12824
rect 16764 12776 16816 12782
rect 16868 12753 16896 15014
rect 16950 14716 17258 14725
rect 16950 14714 16956 14716
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17252 14714 17258 14716
rect 17012 14662 17014 14714
rect 17194 14662 17196 14714
rect 16950 14660 16956 14662
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 17252 14660 17258 14662
rect 16950 14651 17258 14660
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17052 13977 17080 14214
rect 17038 13968 17094 13977
rect 17038 13903 17094 13912
rect 16950 13628 17258 13637
rect 16950 13626 16956 13628
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17252 13626 17258 13628
rect 17012 13574 17014 13626
rect 17194 13574 17196 13626
rect 16950 13572 16956 13574
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 17252 13572 17258 13574
rect 16950 13563 17258 13572
rect 17328 12753 17356 16458
rect 17420 14278 17448 16458
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17512 16153 17540 16390
rect 17610 16348 17918 16357
rect 17610 16346 17616 16348
rect 17672 16346 17696 16348
rect 17752 16346 17776 16348
rect 17832 16346 17856 16348
rect 17912 16346 17918 16348
rect 17672 16294 17674 16346
rect 17854 16294 17856 16346
rect 17610 16292 17616 16294
rect 17672 16292 17696 16294
rect 17752 16292 17776 16294
rect 17832 16292 17856 16294
rect 17912 16292 17918 16294
rect 17610 16283 17918 16292
rect 17498 16144 17554 16153
rect 17498 16079 17554 16088
rect 17972 15910 18000 16390
rect 18156 16114 18184 17614
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 17202 18276 17478
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17972 15558 18276 15586
rect 17972 15366 18000 15558
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17610 15260 17918 15269
rect 17610 15258 17616 15260
rect 17672 15258 17696 15260
rect 17752 15258 17776 15260
rect 17832 15258 17856 15260
rect 17912 15258 17918 15260
rect 17672 15206 17674 15258
rect 17854 15206 17856 15258
rect 17610 15204 17616 15206
rect 17672 15204 17696 15206
rect 17752 15204 17776 15206
rect 17832 15204 17856 15206
rect 17912 15204 17918 15206
rect 17610 15195 17918 15204
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17512 13530 17540 14894
rect 17880 14414 17908 15098
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17610 14172 17918 14181
rect 17610 14170 17616 14172
rect 17672 14170 17696 14172
rect 17752 14170 17776 14172
rect 17832 14170 17856 14172
rect 17912 14170 17918 14172
rect 17672 14118 17674 14170
rect 17854 14118 17856 14170
rect 17610 14116 17616 14118
rect 17672 14116 17696 14118
rect 17752 14116 17776 14118
rect 17832 14116 17856 14118
rect 17912 14116 17918 14118
rect 17610 14107 17918 14116
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17610 13084 17918 13093
rect 17610 13082 17616 13084
rect 17672 13082 17696 13084
rect 17752 13082 17776 13084
rect 17832 13082 17856 13084
rect 17912 13082 17918 13084
rect 17672 13030 17674 13082
rect 17854 13030 17856 13082
rect 17610 13028 17616 13030
rect 17672 13028 17696 13030
rect 17752 13028 17776 13030
rect 17832 13028 17856 13030
rect 17912 13028 17918 13030
rect 17610 13019 17918 13028
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 16764 12718 16816 12724
rect 16854 12744 16910 12753
rect 16776 9722 16804 12718
rect 16854 12679 16910 12688
rect 17314 12744 17370 12753
rect 17314 12679 17370 12688
rect 16950 12540 17258 12549
rect 16950 12538 16956 12540
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17252 12538 17258 12540
rect 17012 12486 17014 12538
rect 17194 12486 17196 12538
rect 16950 12484 16956 12486
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 17252 12484 17258 12486
rect 16950 12475 17258 12484
rect 17406 12336 17462 12345
rect 17406 12271 17462 12280
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 16950 11452 17258 11461
rect 16950 11450 16956 11452
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17252 11450 17258 11452
rect 17012 11398 17014 11450
rect 17194 11398 17196 11450
rect 16950 11396 16956 11398
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 17252 11396 17258 11398
rect 16950 11387 17258 11396
rect 16950 10364 17258 10373
rect 16950 10362 16956 10364
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17252 10362 17258 10364
rect 17012 10310 17014 10362
rect 17194 10310 17196 10362
rect 16950 10308 16956 10310
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 17252 10308 17258 10310
rect 16950 10299 17258 10308
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16868 9602 16896 10066
rect 17040 9988 17092 9994
rect 17040 9930 17092 9936
rect 16776 9586 16988 9602
rect 16776 9580 17000 9586
rect 16776 9574 16948 9580
rect 16776 6798 16804 9574
rect 16948 9522 17000 9528
rect 17052 9466 17080 9930
rect 17132 9512 17184 9518
rect 16868 9438 17080 9466
rect 17130 9480 17132 9489
rect 17184 9480 17186 9489
rect 16868 7546 16896 9438
rect 17130 9415 17186 9424
rect 16950 9276 17258 9285
rect 16950 9274 16956 9276
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17252 9274 17258 9276
rect 17012 9222 17014 9274
rect 17194 9222 17196 9274
rect 16950 9220 16956 9222
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 17252 9220 17258 9222
rect 16950 9211 17258 9220
rect 16950 8188 17258 8197
rect 16950 8186 16956 8188
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17252 8186 17258 8188
rect 17012 8134 17014 8186
rect 17194 8134 17196 8186
rect 16950 8132 16956 8134
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 17252 8132 17258 8134
rect 16950 8123 17258 8132
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16776 5953 16804 6122
rect 16762 5944 16818 5953
rect 16762 5879 16818 5888
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 15660 4616 15712 4622
rect 15658 4584 15660 4593
rect 15712 4584 15714 4593
rect 16316 4554 16344 4762
rect 16776 4622 16804 4966
rect 16868 4826 16896 7346
rect 16950 7100 17258 7109
rect 16950 7098 16956 7100
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17252 7098 17258 7100
rect 17012 7046 17014 7098
rect 17194 7046 17196 7098
rect 16950 7044 16956 7046
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 17252 7044 17258 7046
rect 16950 7035 17258 7044
rect 16950 6012 17258 6021
rect 16950 6010 16956 6012
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17252 6010 17258 6012
rect 17012 5958 17014 6010
rect 17194 5958 17196 6010
rect 16950 5956 16956 5958
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 17252 5956 17258 5958
rect 16950 5947 17258 5956
rect 16950 4924 17258 4933
rect 16950 4922 16956 4924
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17252 4922 17258 4924
rect 17012 4870 17014 4922
rect 17194 4870 17196 4922
rect 16950 4868 16956 4870
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 17252 4868 17258 4870
rect 16950 4859 17258 4868
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 15658 4519 15714 4528
rect 16304 4548 16356 4554
rect 16304 4490 16356 4496
rect 16396 4548 16448 4554
rect 16396 4490 16448 4496
rect 16408 4214 16436 4490
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15750 2544 15806 2553
rect 15750 2479 15806 2488
rect 15764 2446 15792 2479
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 16118 2408 16174 2417
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 13728 2372 13780 2378
rect 16224 2378 16252 3878
rect 16950 3836 17258 3845
rect 16950 3834 16956 3836
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17252 3834 17258 3836
rect 17012 3782 17014 3834
rect 17194 3782 17196 3834
rect 16950 3780 16956 3782
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 17252 3780 17258 3782
rect 16950 3771 17258 3780
rect 17328 3738 17356 11630
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 16950 2748 17258 2757
rect 16950 2746 16956 2748
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17252 2746 17258 2748
rect 17012 2694 17014 2746
rect 17194 2694 17196 2746
rect 16950 2692 16956 2694
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 17252 2692 17258 2694
rect 16950 2683 17258 2692
rect 17420 2582 17448 12271
rect 17512 9042 17540 12854
rect 17610 11996 17918 12005
rect 17610 11994 17616 11996
rect 17672 11994 17696 11996
rect 17752 11994 17776 11996
rect 17832 11994 17856 11996
rect 17912 11994 17918 11996
rect 17672 11942 17674 11994
rect 17854 11942 17856 11994
rect 17610 11940 17616 11942
rect 17672 11940 17696 11942
rect 17752 11940 17776 11942
rect 17832 11940 17856 11942
rect 17912 11940 17918 11942
rect 17610 11931 17918 11940
rect 17610 10908 17918 10917
rect 17610 10906 17616 10908
rect 17672 10906 17696 10908
rect 17752 10906 17776 10908
rect 17832 10906 17856 10908
rect 17912 10906 17918 10908
rect 17672 10854 17674 10906
rect 17854 10854 17856 10906
rect 17610 10852 17616 10854
rect 17672 10852 17696 10854
rect 17752 10852 17776 10854
rect 17832 10852 17856 10854
rect 17912 10852 17918 10854
rect 17610 10843 17918 10852
rect 17972 10538 18000 15030
rect 18064 12238 18092 15438
rect 18156 13734 18184 15438
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 10266 17816 10406
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17972 10198 18000 10474
rect 17960 10192 18012 10198
rect 17866 10160 17922 10169
rect 17960 10134 18012 10140
rect 17866 10095 17868 10104
rect 17920 10095 17922 10104
rect 17868 10066 17920 10072
rect 17610 9820 17918 9829
rect 17610 9818 17616 9820
rect 17672 9818 17696 9820
rect 17752 9818 17776 9820
rect 17832 9818 17856 9820
rect 17912 9818 17918 9820
rect 17672 9766 17674 9818
rect 17854 9766 17856 9818
rect 17610 9764 17616 9766
rect 17672 9764 17696 9766
rect 17752 9764 17776 9766
rect 17832 9764 17856 9766
rect 17912 9764 17918 9766
rect 17610 9755 17918 9764
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17512 8090 17540 8842
rect 17604 8838 17632 9318
rect 17592 8832 17644 8838
rect 17880 8820 17908 9454
rect 18064 9178 18092 12174
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17958 9072 18014 9081
rect 17958 9007 18014 9016
rect 17972 8974 18000 9007
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17880 8792 18000 8820
rect 17592 8774 17644 8780
rect 17610 8732 17918 8741
rect 17610 8730 17616 8732
rect 17672 8730 17696 8732
rect 17752 8730 17776 8732
rect 17832 8730 17856 8732
rect 17912 8730 17918 8732
rect 17672 8678 17674 8730
rect 17854 8678 17856 8730
rect 17610 8676 17616 8678
rect 17672 8676 17696 8678
rect 17752 8676 17776 8678
rect 17832 8676 17856 8678
rect 17912 8676 17918 8678
rect 17610 8667 17918 8676
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17682 7984 17738 7993
rect 17682 7919 17738 7928
rect 17696 7886 17724 7919
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17610 7644 17918 7653
rect 17610 7642 17616 7644
rect 17672 7642 17696 7644
rect 17752 7642 17776 7644
rect 17832 7642 17856 7644
rect 17912 7642 17918 7644
rect 17672 7590 17674 7642
rect 17854 7590 17856 7642
rect 17610 7588 17616 7590
rect 17672 7588 17696 7590
rect 17752 7588 17776 7590
rect 17832 7588 17856 7590
rect 17912 7588 17918 7590
rect 17610 7579 17918 7588
rect 17610 6556 17918 6565
rect 17610 6554 17616 6556
rect 17672 6554 17696 6556
rect 17752 6554 17776 6556
rect 17832 6554 17856 6556
rect 17912 6554 17918 6556
rect 17672 6502 17674 6554
rect 17854 6502 17856 6554
rect 17610 6500 17616 6502
rect 17672 6500 17696 6502
rect 17752 6500 17776 6502
rect 17832 6500 17856 6502
rect 17912 6500 17918 6502
rect 17610 6491 17918 6500
rect 17610 5468 17918 5477
rect 17610 5466 17616 5468
rect 17672 5466 17696 5468
rect 17752 5466 17776 5468
rect 17832 5466 17856 5468
rect 17912 5466 17918 5468
rect 17672 5414 17674 5466
rect 17854 5414 17856 5466
rect 17610 5412 17616 5414
rect 17672 5412 17696 5414
rect 17752 5412 17776 5414
rect 17832 5412 17856 5414
rect 17912 5412 17918 5414
rect 17610 5403 17918 5412
rect 17610 4380 17918 4389
rect 17610 4378 17616 4380
rect 17672 4378 17696 4380
rect 17752 4378 17776 4380
rect 17832 4378 17856 4380
rect 17912 4378 17918 4380
rect 17672 4326 17674 4378
rect 17854 4326 17856 4378
rect 17610 4324 17616 4326
rect 17672 4324 17696 4326
rect 17752 4324 17776 4326
rect 17832 4324 17856 4326
rect 17912 4324 17918 4326
rect 17610 4315 17918 4324
rect 17972 4214 18000 8792
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17512 2514 17540 4150
rect 17610 3292 17918 3301
rect 17610 3290 17616 3292
rect 17672 3290 17696 3292
rect 17752 3290 17776 3292
rect 17832 3290 17856 3292
rect 17912 3290 17918 3292
rect 17672 3238 17674 3290
rect 17854 3238 17856 3290
rect 17610 3236 17616 3238
rect 17672 3236 17696 3238
rect 17752 3236 17776 3238
rect 17832 3236 17856 3238
rect 17912 3236 17918 3238
rect 17610 3227 17918 3236
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 16118 2343 16120 2352
rect 13728 2314 13780 2320
rect 16172 2343 16174 2352
rect 16212 2372 16264 2378
rect 16120 2314 16172 2320
rect 16212 2314 16264 2320
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 1858 1728 1914 1737
rect 1858 1663 1914 1672
rect 3344 800 3372 2314
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 9968 800 9996 2314
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 16592 800 16620 2382
rect 18064 2378 18092 8570
rect 18156 6458 18184 11630
rect 18248 10062 18276 15558
rect 18340 15162 18368 16730
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18340 9586 18368 14962
rect 18432 14482 18460 16390
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18432 13705 18460 14010
rect 18418 13696 18474 13705
rect 18418 13631 18474 13640
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11257 18460 11494
rect 18418 11248 18474 11257
rect 18418 11183 18474 11192
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18432 9926 18460 10406
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18248 6474 18276 9454
rect 18432 9450 18460 9862
rect 18420 9444 18472 9450
rect 18420 9386 18472 9392
rect 18420 8832 18472 8838
rect 18418 8800 18420 8809
rect 18472 8800 18474 8809
rect 18418 8735 18474 8744
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18144 6452 18196 6458
rect 18248 6446 18368 6474
rect 18144 6394 18196 6400
rect 18234 6352 18290 6361
rect 18234 6287 18290 6296
rect 18248 6254 18276 6287
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18340 6118 18368 6446
rect 18432 6361 18460 6598
rect 18418 6352 18474 6361
rect 18418 6287 18474 6296
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 18236 5636 18288 5642
rect 18236 5578 18288 5584
rect 18248 4146 18276 5578
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18340 4078 18368 6054
rect 18524 4758 18552 16662
rect 18788 16652 18840 16658
rect 18788 16594 18840 16600
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18616 15026 18644 16050
rect 18696 15428 18748 15434
rect 18696 15370 18748 15376
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18708 11898 18736 15370
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18604 11620 18656 11626
rect 18604 11562 18656 11568
rect 18512 4752 18564 4758
rect 18512 4694 18564 4700
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18420 3936 18472 3942
rect 18418 3904 18420 3913
rect 18472 3904 18474 3913
rect 18418 3839 18474 3848
rect 18616 2446 18644 11562
rect 18708 2854 18736 11698
rect 18800 6798 18828 16594
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18892 14822 18920 16118
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18892 9042 18920 14758
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18984 7750 19012 11834
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 17610 2204 17918 2213
rect 17610 2202 17616 2204
rect 17672 2202 17696 2204
rect 17752 2202 17776 2204
rect 17832 2202 17856 2204
rect 17912 2202 17918 2204
rect 17672 2150 17674 2202
rect 17854 2150 17856 2202
rect 17610 2148 17616 2150
rect 17672 2148 17696 2150
rect 17752 2148 17776 2150
rect 17832 2148 17856 2150
rect 17912 2148 17918 2150
rect 17610 2139 17918 2148
rect 18432 1465 18460 2246
rect 18418 1456 18474 1465
rect 18418 1391 18474 1400
rect 3330 0 3386 800
rect 9954 0 10010 800
rect 16578 0 16634 800
<< via2 >>
rect 17866 18536 17922 18592
rect 1858 17992 1914 18048
rect 2616 17434 2672 17436
rect 2696 17434 2752 17436
rect 2776 17434 2832 17436
rect 2856 17434 2912 17436
rect 2616 17382 2662 17434
rect 2662 17382 2672 17434
rect 2696 17382 2726 17434
rect 2726 17382 2738 17434
rect 2738 17382 2752 17434
rect 2776 17382 2790 17434
rect 2790 17382 2802 17434
rect 2802 17382 2832 17434
rect 2856 17382 2866 17434
rect 2866 17382 2912 17434
rect 2616 17380 2672 17382
rect 2696 17380 2752 17382
rect 2776 17380 2832 17382
rect 2856 17380 2912 17382
rect 846 17040 902 17096
rect 1030 15816 1086 15872
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 1490 15972 1546 16008
rect 1490 15952 1492 15972
rect 1492 15952 1544 15972
rect 1544 15952 1546 15972
rect 846 14864 902 14920
rect 1398 13640 1454 13696
rect 846 12688 902 12744
rect 846 11600 902 11656
rect 1306 11192 1362 11248
rect 1214 10648 1270 10704
rect 846 10240 902 10296
rect 846 9424 902 9480
rect 846 7248 902 7304
rect 938 6024 994 6080
rect 846 5072 902 5128
rect 846 3984 902 4040
rect 846 2896 902 2952
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 1398 9968 1454 10024
rect 1398 8200 1454 8256
rect 2616 16346 2672 16348
rect 2696 16346 2752 16348
rect 2776 16346 2832 16348
rect 2856 16346 2912 16348
rect 2616 16294 2662 16346
rect 2662 16294 2672 16346
rect 2696 16294 2726 16346
rect 2726 16294 2738 16346
rect 2738 16294 2752 16346
rect 2776 16294 2790 16346
rect 2790 16294 2802 16346
rect 2802 16294 2832 16346
rect 2856 16294 2866 16346
rect 2866 16294 2912 16346
rect 2616 16292 2672 16294
rect 2696 16292 2752 16294
rect 2776 16292 2832 16294
rect 2856 16292 2912 16294
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 1766 6180 1822 6216
rect 1766 6160 1768 6180
rect 1768 6160 1820 6180
rect 1820 6160 1822 6180
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 3054 15952 3110 16008
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 2502 9968 2558 10024
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 2594 8880 2650 8936
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 2318 7828 2320 7848
rect 2320 7828 2372 7848
rect 2372 7828 2374 7848
rect 2318 7792 2374 7828
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 2042 6704 2098 6760
rect 3514 13776 3570 13832
rect 3146 9716 3202 9752
rect 3146 9696 3148 9716
rect 3148 9696 3200 9716
rect 3200 9696 3202 9716
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 4710 16360 4766 16416
rect 3790 10784 3846 10840
rect 3698 9424 3754 9480
rect 3974 15000 4030 15056
rect 4342 15544 4398 15600
rect 3974 11600 4030 11656
rect 3422 8336 3478 8392
rect 3146 5208 3202 5264
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 4066 8880 4122 8936
rect 4066 8744 4122 8800
rect 4434 12844 4490 12880
rect 4434 12824 4436 12844
rect 4436 12824 4488 12844
rect 4488 12824 4490 12844
rect 4802 15988 4804 16008
rect 4804 15988 4856 16008
rect 4856 15988 4858 16008
rect 4802 15952 4858 15988
rect 4894 13368 4950 13424
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 2318 2896 2374 2952
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 7616 17434 7672 17436
rect 7696 17434 7752 17436
rect 7776 17434 7832 17436
rect 7856 17434 7912 17436
rect 7616 17382 7662 17434
rect 7662 17382 7672 17434
rect 7696 17382 7726 17434
rect 7726 17382 7738 17434
rect 7738 17382 7752 17434
rect 7776 17382 7790 17434
rect 7790 17382 7802 17434
rect 7802 17382 7832 17434
rect 7856 17382 7866 17434
rect 7866 17382 7912 17434
rect 7616 17380 7672 17382
rect 7696 17380 7752 17382
rect 7776 17380 7832 17382
rect 7856 17380 7912 17382
rect 6956 16890 7012 16892
rect 7036 16890 7092 16892
rect 7116 16890 7172 16892
rect 7196 16890 7252 16892
rect 6956 16838 7002 16890
rect 7002 16838 7012 16890
rect 7036 16838 7066 16890
rect 7066 16838 7078 16890
rect 7078 16838 7092 16890
rect 7116 16838 7130 16890
rect 7130 16838 7142 16890
rect 7142 16838 7172 16890
rect 7196 16838 7206 16890
rect 7206 16838 7252 16890
rect 6956 16836 7012 16838
rect 7036 16836 7092 16838
rect 7116 16836 7172 16838
rect 7196 16836 7252 16838
rect 5354 15952 5410 16008
rect 5354 11328 5410 11384
rect 5078 10140 5080 10160
rect 5080 10140 5132 10160
rect 5132 10140 5134 10160
rect 5078 10104 5134 10140
rect 5538 9968 5594 10024
rect 4894 6704 4950 6760
rect 6090 10512 6146 10568
rect 5170 5092 5226 5128
rect 5170 5072 5172 5092
rect 5172 5072 5224 5092
rect 5224 5072 5226 5092
rect 6642 15272 6698 15328
rect 6918 16496 6974 16552
rect 6956 15802 7012 15804
rect 7036 15802 7092 15804
rect 7116 15802 7172 15804
rect 7196 15802 7252 15804
rect 6956 15750 7002 15802
rect 7002 15750 7012 15802
rect 7036 15750 7066 15802
rect 7066 15750 7078 15802
rect 7078 15750 7092 15802
rect 7116 15750 7130 15802
rect 7130 15750 7142 15802
rect 7142 15750 7172 15802
rect 7196 15750 7206 15802
rect 7206 15750 7252 15802
rect 6956 15748 7012 15750
rect 7036 15748 7092 15750
rect 7116 15748 7172 15750
rect 7196 15748 7252 15750
rect 6458 11056 6514 11112
rect 6956 14714 7012 14716
rect 7036 14714 7092 14716
rect 7116 14714 7172 14716
rect 7196 14714 7252 14716
rect 6956 14662 7002 14714
rect 7002 14662 7012 14714
rect 7036 14662 7066 14714
rect 7066 14662 7078 14714
rect 7078 14662 7092 14714
rect 7116 14662 7130 14714
rect 7130 14662 7142 14714
rect 7142 14662 7172 14714
rect 7196 14662 7206 14714
rect 7206 14662 7252 14714
rect 6956 14660 7012 14662
rect 7036 14660 7092 14662
rect 7116 14660 7172 14662
rect 7196 14660 7252 14662
rect 6826 14456 6882 14512
rect 6734 11328 6790 11384
rect 6550 9016 6606 9072
rect 6458 8744 6514 8800
rect 6274 4120 6330 4176
rect 5814 4004 5870 4040
rect 5814 3984 5816 4004
rect 5816 3984 5868 4004
rect 5868 3984 5870 4004
rect 6642 8372 6644 8392
rect 6644 8372 6696 8392
rect 6696 8372 6698 8392
rect 6642 8336 6698 8372
rect 6956 13626 7012 13628
rect 7036 13626 7092 13628
rect 7116 13626 7172 13628
rect 7196 13626 7252 13628
rect 6956 13574 7002 13626
rect 7002 13574 7012 13626
rect 7036 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7092 13626
rect 7116 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7172 13626
rect 7196 13574 7206 13626
rect 7206 13574 7252 13626
rect 6956 13572 7012 13574
rect 7036 13572 7092 13574
rect 7116 13572 7172 13574
rect 7196 13572 7252 13574
rect 7010 12688 7066 12744
rect 7194 12688 7250 12744
rect 7470 16360 7526 16416
rect 8022 16360 8078 16416
rect 7616 16346 7672 16348
rect 7696 16346 7752 16348
rect 7776 16346 7832 16348
rect 7856 16346 7912 16348
rect 7616 16294 7662 16346
rect 7662 16294 7672 16346
rect 7696 16294 7726 16346
rect 7726 16294 7738 16346
rect 7738 16294 7752 16346
rect 7776 16294 7790 16346
rect 7790 16294 7802 16346
rect 7802 16294 7832 16346
rect 7856 16294 7866 16346
rect 7866 16294 7912 16346
rect 7616 16292 7672 16294
rect 7696 16292 7752 16294
rect 7776 16292 7832 16294
rect 7856 16292 7912 16294
rect 7616 15258 7672 15260
rect 7696 15258 7752 15260
rect 7776 15258 7832 15260
rect 7856 15258 7912 15260
rect 7616 15206 7662 15258
rect 7662 15206 7672 15258
rect 7696 15206 7726 15258
rect 7726 15206 7738 15258
rect 7738 15206 7752 15258
rect 7776 15206 7790 15258
rect 7790 15206 7802 15258
rect 7802 15206 7832 15258
rect 7856 15206 7866 15258
rect 7866 15206 7912 15258
rect 7616 15204 7672 15206
rect 7696 15204 7752 15206
rect 7776 15204 7832 15206
rect 7856 15204 7912 15206
rect 7616 14170 7672 14172
rect 7696 14170 7752 14172
rect 7776 14170 7832 14172
rect 7856 14170 7912 14172
rect 7616 14118 7662 14170
rect 7662 14118 7672 14170
rect 7696 14118 7726 14170
rect 7726 14118 7738 14170
rect 7738 14118 7752 14170
rect 7776 14118 7790 14170
rect 7790 14118 7802 14170
rect 7802 14118 7832 14170
rect 7856 14118 7866 14170
rect 7866 14118 7912 14170
rect 7616 14116 7672 14118
rect 7696 14116 7752 14118
rect 7776 14116 7832 14118
rect 7856 14116 7912 14118
rect 7562 13232 7618 13288
rect 7616 13082 7672 13084
rect 7696 13082 7752 13084
rect 7776 13082 7832 13084
rect 7856 13082 7912 13084
rect 7616 13030 7662 13082
rect 7662 13030 7672 13082
rect 7696 13030 7726 13082
rect 7726 13030 7738 13082
rect 7738 13030 7752 13082
rect 7776 13030 7790 13082
rect 7790 13030 7802 13082
rect 7802 13030 7832 13082
rect 7856 13030 7866 13082
rect 7866 13030 7912 13082
rect 7616 13028 7672 13030
rect 7696 13028 7752 13030
rect 7776 13028 7832 13030
rect 7856 13028 7912 13030
rect 6956 12538 7012 12540
rect 7036 12538 7092 12540
rect 7116 12538 7172 12540
rect 7196 12538 7252 12540
rect 6956 12486 7002 12538
rect 7002 12486 7012 12538
rect 7036 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7092 12538
rect 7116 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7172 12538
rect 7196 12486 7206 12538
rect 7206 12486 7252 12538
rect 6956 12484 7012 12486
rect 7036 12484 7092 12486
rect 7116 12484 7172 12486
rect 7196 12484 7252 12486
rect 7194 12164 7250 12200
rect 7194 12144 7196 12164
rect 7196 12144 7248 12164
rect 7248 12144 7250 12164
rect 7286 11756 7342 11792
rect 7286 11736 7288 11756
rect 7288 11736 7340 11756
rect 7340 11736 7342 11756
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 7286 9716 7342 9752
rect 7286 9696 7288 9716
rect 7288 9696 7340 9716
rect 7340 9696 7342 9716
rect 6918 9424 6974 9480
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 7746 12588 7748 12608
rect 7748 12588 7800 12608
rect 7800 12588 7802 12608
rect 7746 12552 7802 12588
rect 7746 12280 7802 12336
rect 8298 13368 8354 13424
rect 8390 12552 8446 12608
rect 8390 12280 8446 12336
rect 8298 12144 8354 12200
rect 7616 11994 7672 11996
rect 7696 11994 7752 11996
rect 7776 11994 7832 11996
rect 7856 11994 7912 11996
rect 7616 11942 7662 11994
rect 7662 11942 7672 11994
rect 7696 11942 7726 11994
rect 7726 11942 7738 11994
rect 7738 11942 7752 11994
rect 7776 11942 7790 11994
rect 7790 11942 7802 11994
rect 7802 11942 7832 11994
rect 7856 11942 7866 11994
rect 7866 11942 7912 11994
rect 7616 11940 7672 11942
rect 7696 11940 7752 11942
rect 7776 11940 7832 11942
rect 7856 11940 7912 11942
rect 7838 11600 7894 11656
rect 8022 11600 8078 11656
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 7562 10240 7618 10296
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 6734 5752 6790 5808
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 7654 8336 7710 8392
rect 7378 8200 7434 8256
rect 7930 7792 7986 7848
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 8666 13812 8668 13832
rect 8668 13812 8720 13832
rect 8720 13812 8722 13832
rect 8666 13776 8722 13812
rect 8666 12824 8722 12880
rect 9034 15544 9090 15600
rect 9126 15408 9182 15464
rect 9126 13776 9182 13832
rect 8850 12688 8906 12744
rect 8114 8064 8170 8120
rect 8298 9832 8354 9888
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 8666 6704 8722 6760
rect 12616 17434 12672 17436
rect 12696 17434 12752 17436
rect 12776 17434 12832 17436
rect 12856 17434 12912 17436
rect 12616 17382 12662 17434
rect 12662 17382 12672 17434
rect 12696 17382 12726 17434
rect 12726 17382 12738 17434
rect 12738 17382 12752 17434
rect 12776 17382 12790 17434
rect 12790 17382 12802 17434
rect 12802 17382 12832 17434
rect 12856 17382 12866 17434
rect 12866 17382 12912 17434
rect 12616 17380 12672 17382
rect 12696 17380 12752 17382
rect 12776 17380 12832 17382
rect 12856 17380 12912 17382
rect 9402 16224 9458 16280
rect 9402 15272 9458 15328
rect 8942 8744 8998 8800
rect 8942 5072 8998 5128
rect 8850 3576 8906 3632
rect 9034 4392 9090 4448
rect 9770 15408 9826 15464
rect 9678 15156 9734 15192
rect 9678 15136 9680 15156
rect 9680 15136 9732 15156
rect 9732 15136 9734 15156
rect 9770 14900 9772 14920
rect 9772 14900 9824 14920
rect 9824 14900 9826 14920
rect 9770 14864 9826 14900
rect 9678 14728 9734 14784
rect 9678 14612 9734 14648
rect 9678 14592 9680 14612
rect 9680 14592 9732 14612
rect 9732 14592 9734 14612
rect 9586 14320 9642 14376
rect 9770 14456 9826 14512
rect 9586 13252 9642 13288
rect 9586 13232 9588 13252
rect 9588 13232 9640 13252
rect 9640 13232 9642 13252
rect 9494 12416 9550 12472
rect 9678 12688 9734 12744
rect 9678 12300 9734 12336
rect 9678 12280 9680 12300
rect 9680 12280 9732 12300
rect 9732 12280 9734 12300
rect 9494 11736 9550 11792
rect 9586 9560 9642 9616
rect 9862 12824 9918 12880
rect 9770 10104 9826 10160
rect 9770 8336 9826 8392
rect 10046 15680 10102 15736
rect 10138 15000 10194 15056
rect 10322 16532 10324 16552
rect 10324 16532 10376 16552
rect 10376 16532 10378 16552
rect 10322 16496 10378 16532
rect 10414 15272 10470 15328
rect 10322 15136 10378 15192
rect 10690 15408 10746 15464
rect 10598 15272 10654 15328
rect 10138 13912 10194 13968
rect 10322 13912 10378 13968
rect 10598 14728 10654 14784
rect 10506 14592 10562 14648
rect 10598 14456 10654 14512
rect 10322 9696 10378 9752
rect 9954 4256 10010 4312
rect 10138 3984 10194 4040
rect 10506 11872 10562 11928
rect 10966 15272 11022 15328
rect 10966 15136 11022 15192
rect 11058 12552 11114 12608
rect 9126 2624 9182 2680
rect 11242 12552 11298 12608
rect 11150 4800 11206 4856
rect 10966 3188 11022 3224
rect 10966 3168 10968 3188
rect 10968 3168 11020 3188
rect 11020 3168 11022 3188
rect 11426 15408 11482 15464
rect 11426 14184 11482 14240
rect 11956 16890 12012 16892
rect 12036 16890 12092 16892
rect 12116 16890 12172 16892
rect 12196 16890 12252 16892
rect 11956 16838 12002 16890
rect 12002 16838 12012 16890
rect 12036 16838 12066 16890
rect 12066 16838 12078 16890
rect 12078 16838 12092 16890
rect 12116 16838 12130 16890
rect 12130 16838 12142 16890
rect 12142 16838 12172 16890
rect 12196 16838 12206 16890
rect 12206 16838 12252 16890
rect 11956 16836 12012 16838
rect 12036 16836 12092 16838
rect 12116 16836 12172 16838
rect 12196 16836 12252 16838
rect 11978 16224 12034 16280
rect 12254 16088 12310 16144
rect 11956 15802 12012 15804
rect 12036 15802 12092 15804
rect 12116 15802 12172 15804
rect 12196 15802 12252 15804
rect 11956 15750 12002 15802
rect 12002 15750 12012 15802
rect 12036 15750 12066 15802
rect 12066 15750 12078 15802
rect 12078 15750 12092 15802
rect 12116 15750 12130 15802
rect 12130 15750 12142 15802
rect 12142 15750 12172 15802
rect 12196 15750 12206 15802
rect 12206 15750 12252 15802
rect 11956 15748 12012 15750
rect 12036 15748 12092 15750
rect 12116 15748 12172 15750
rect 12196 15748 12252 15750
rect 12346 14728 12402 14784
rect 11956 14714 12012 14716
rect 12036 14714 12092 14716
rect 12116 14714 12172 14716
rect 12196 14714 12252 14716
rect 11956 14662 12002 14714
rect 12002 14662 12012 14714
rect 12036 14662 12066 14714
rect 12066 14662 12078 14714
rect 12078 14662 12092 14714
rect 12116 14662 12130 14714
rect 12130 14662 12142 14714
rect 12142 14662 12172 14714
rect 12196 14662 12206 14714
rect 12206 14662 12252 14714
rect 11956 14660 12012 14662
rect 12036 14660 12092 14662
rect 12116 14660 12172 14662
rect 12196 14660 12252 14662
rect 11956 13626 12012 13628
rect 12036 13626 12092 13628
rect 12116 13626 12172 13628
rect 12196 13626 12252 13628
rect 11956 13574 12002 13626
rect 12002 13574 12012 13626
rect 12036 13574 12066 13626
rect 12066 13574 12078 13626
rect 12078 13574 12092 13626
rect 12116 13574 12130 13626
rect 12130 13574 12142 13626
rect 12142 13574 12172 13626
rect 12196 13574 12206 13626
rect 12206 13574 12252 13626
rect 11956 13572 12012 13574
rect 12036 13572 12092 13574
rect 12116 13572 12172 13574
rect 12196 13572 12252 13574
rect 11702 12280 11758 12336
rect 11518 11328 11574 11384
rect 11956 12538 12012 12540
rect 12036 12538 12092 12540
rect 12116 12538 12172 12540
rect 12196 12538 12252 12540
rect 11956 12486 12002 12538
rect 12002 12486 12012 12538
rect 12036 12486 12066 12538
rect 12066 12486 12078 12538
rect 12078 12486 12092 12538
rect 12116 12486 12130 12538
rect 12130 12486 12142 12538
rect 12142 12486 12172 12538
rect 12196 12486 12206 12538
rect 12206 12486 12252 12538
rect 11956 12484 12012 12486
rect 12036 12484 12092 12486
rect 12116 12484 12172 12486
rect 12196 12484 12252 12486
rect 11978 12280 12034 12336
rect 11886 11872 11942 11928
rect 11956 11450 12012 11452
rect 12036 11450 12092 11452
rect 12116 11450 12172 11452
rect 12196 11450 12252 11452
rect 11956 11398 12002 11450
rect 12002 11398 12012 11450
rect 12036 11398 12066 11450
rect 12066 11398 12078 11450
rect 12078 11398 12092 11450
rect 12116 11398 12130 11450
rect 12130 11398 12142 11450
rect 12142 11398 12172 11450
rect 12196 11398 12206 11450
rect 12206 11398 12252 11450
rect 11956 11396 12012 11398
rect 12036 11396 12092 11398
rect 12116 11396 12172 11398
rect 12196 11396 12252 11398
rect 11794 10784 11850 10840
rect 11702 9424 11758 9480
rect 11702 8744 11758 8800
rect 11956 10362 12012 10364
rect 12036 10362 12092 10364
rect 12116 10362 12172 10364
rect 12196 10362 12252 10364
rect 11956 10310 12002 10362
rect 12002 10310 12012 10362
rect 12036 10310 12066 10362
rect 12066 10310 12078 10362
rect 12078 10310 12092 10362
rect 12116 10310 12130 10362
rect 12130 10310 12142 10362
rect 12142 10310 12172 10362
rect 12196 10310 12206 10362
rect 12206 10310 12252 10362
rect 11956 10308 12012 10310
rect 12036 10308 12092 10310
rect 12116 10308 12172 10310
rect 12196 10308 12252 10310
rect 11956 9274 12012 9276
rect 12036 9274 12092 9276
rect 12116 9274 12172 9276
rect 12196 9274 12252 9276
rect 11956 9222 12002 9274
rect 12002 9222 12012 9274
rect 12036 9222 12066 9274
rect 12066 9222 12078 9274
rect 12078 9222 12092 9274
rect 12116 9222 12130 9274
rect 12130 9222 12142 9274
rect 12142 9222 12172 9274
rect 12196 9222 12206 9274
rect 12206 9222 12252 9274
rect 11956 9220 12012 9222
rect 12036 9220 12092 9222
rect 12116 9220 12172 9222
rect 12196 9220 12252 9222
rect 13266 16360 13322 16416
rect 12616 16346 12672 16348
rect 12696 16346 12752 16348
rect 12776 16346 12832 16348
rect 12856 16346 12912 16348
rect 12616 16294 12662 16346
rect 12662 16294 12672 16346
rect 12696 16294 12726 16346
rect 12726 16294 12738 16346
rect 12738 16294 12752 16346
rect 12776 16294 12790 16346
rect 12790 16294 12802 16346
rect 12802 16294 12832 16346
rect 12856 16294 12866 16346
rect 12866 16294 12912 16346
rect 12616 16292 12672 16294
rect 12696 16292 12752 16294
rect 12776 16292 12832 16294
rect 12856 16292 12912 16294
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 12530 14592 12586 14648
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 12990 13640 13046 13696
rect 12714 13368 12770 13424
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 13634 15952 13690 16008
rect 13542 15564 13598 15600
rect 13542 15544 13544 15564
rect 13544 15544 13596 15564
rect 13596 15544 13598 15564
rect 14094 17040 14150 17096
rect 13634 13812 13636 13832
rect 13636 13812 13688 13832
rect 13688 13812 13690 13832
rect 13634 13776 13690 13812
rect 13450 13640 13506 13696
rect 13082 12980 13138 13016
rect 13082 12960 13084 12980
rect 13084 12960 13136 12980
rect 13136 12960 13138 12980
rect 12622 12416 12678 12472
rect 12990 12316 12992 12336
rect 12992 12316 13044 12336
rect 13044 12316 13046 12336
rect 12990 12280 13046 12316
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 13266 12280 13322 12336
rect 12990 11600 13046 11656
rect 12714 11464 12770 11520
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 11956 8186 12012 8188
rect 12036 8186 12092 8188
rect 12116 8186 12172 8188
rect 12196 8186 12252 8188
rect 11956 8134 12002 8186
rect 12002 8134 12012 8186
rect 12036 8134 12066 8186
rect 12066 8134 12078 8186
rect 12078 8134 12092 8186
rect 12116 8134 12130 8186
rect 12130 8134 12142 8186
rect 12142 8134 12172 8186
rect 12196 8134 12206 8186
rect 12206 8134 12252 8186
rect 11956 8132 12012 8134
rect 12036 8132 12092 8134
rect 12116 8132 12172 8134
rect 12196 8132 12252 8134
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 11956 7098 12012 7100
rect 12036 7098 12092 7100
rect 12116 7098 12172 7100
rect 12196 7098 12252 7100
rect 11956 7046 12002 7098
rect 12002 7046 12012 7098
rect 12036 7046 12066 7098
rect 12066 7046 12078 7098
rect 12078 7046 12092 7098
rect 12116 7046 12130 7098
rect 12130 7046 12142 7098
rect 12142 7046 12172 7098
rect 12196 7046 12206 7098
rect 12206 7046 12252 7098
rect 11956 7044 12012 7046
rect 12036 7044 12092 7046
rect 12116 7044 12172 7046
rect 12196 7044 12252 7046
rect 12530 6840 12586 6896
rect 11956 6010 12012 6012
rect 12036 6010 12092 6012
rect 12116 6010 12172 6012
rect 12196 6010 12252 6012
rect 11956 5958 12002 6010
rect 12002 5958 12012 6010
rect 12036 5958 12066 6010
rect 12066 5958 12078 6010
rect 12078 5958 12092 6010
rect 12116 5958 12130 6010
rect 12130 5958 12142 6010
rect 12142 5958 12172 6010
rect 12196 5958 12206 6010
rect 12206 5958 12252 6010
rect 11956 5956 12012 5958
rect 12036 5956 12092 5958
rect 12116 5956 12172 5958
rect 12196 5956 12252 5958
rect 12254 5228 12310 5264
rect 12254 5208 12256 5228
rect 12256 5208 12308 5228
rect 12308 5208 12310 5228
rect 11956 4922 12012 4924
rect 12036 4922 12092 4924
rect 12116 4922 12172 4924
rect 12196 4922 12252 4924
rect 11956 4870 12002 4922
rect 12002 4870 12012 4922
rect 12036 4870 12066 4922
rect 12066 4870 12078 4922
rect 12078 4870 12092 4922
rect 12116 4870 12130 4922
rect 12130 4870 12142 4922
rect 12142 4870 12172 4922
rect 12196 4870 12206 4922
rect 12206 4870 12252 4922
rect 11956 4868 12012 4870
rect 12036 4868 12092 4870
rect 12116 4868 12172 4870
rect 12196 4868 12252 4870
rect 12070 4700 12072 4720
rect 12072 4700 12124 4720
rect 12124 4700 12126 4720
rect 12070 4664 12126 4700
rect 12254 4664 12310 4720
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 13266 8880 13322 8936
rect 13818 13812 13820 13832
rect 13820 13812 13872 13832
rect 13872 13812 13874 13832
rect 13818 13776 13874 13812
rect 13450 12416 13506 12472
rect 13450 12044 13452 12064
rect 13452 12044 13504 12064
rect 13504 12044 13506 12064
rect 13450 12008 13506 12044
rect 14186 16516 14242 16552
rect 14186 16496 14188 16516
rect 14188 16496 14240 16516
rect 14240 16496 14242 16516
rect 14002 12824 14058 12880
rect 13818 10668 13874 10704
rect 13818 10648 13820 10668
rect 13820 10648 13872 10668
rect 13872 10648 13874 10668
rect 15198 16632 15254 16688
rect 14370 14900 14372 14920
rect 14372 14900 14424 14920
rect 14424 14900 14426 14920
rect 14370 14864 14426 14900
rect 14278 14592 14334 14648
rect 14554 14456 14610 14512
rect 14554 13268 14556 13288
rect 14556 13268 14608 13288
rect 14608 13268 14610 13288
rect 14554 13232 14610 13268
rect 14186 11328 14242 11384
rect 13818 6840 13874 6896
rect 13726 6432 13782 6488
rect 13818 5888 13874 5944
rect 13174 5108 13176 5128
rect 13176 5108 13228 5128
rect 13228 5108 13230 5128
rect 13174 5072 13230 5108
rect 12346 4392 12402 4448
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 12254 4120 12310 4176
rect 12346 4004 12402 4040
rect 12346 3984 12348 4004
rect 12348 3984 12400 4004
rect 12400 3984 12402 4004
rect 11956 3834 12012 3836
rect 12036 3834 12092 3836
rect 12116 3834 12172 3836
rect 12196 3834 12252 3836
rect 11956 3782 12002 3834
rect 12002 3782 12012 3834
rect 12036 3782 12066 3834
rect 12066 3782 12078 3834
rect 12078 3782 12092 3834
rect 12116 3782 12130 3834
rect 12130 3782 12142 3834
rect 12142 3782 12172 3834
rect 12196 3782 12206 3834
rect 12206 3782 12252 3834
rect 11956 3780 12012 3782
rect 12036 3780 12092 3782
rect 12116 3780 12172 3782
rect 12196 3780 12252 3782
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 11956 2746 12012 2748
rect 12036 2746 12092 2748
rect 12116 2746 12172 2748
rect 12196 2746 12252 2748
rect 11956 2694 12002 2746
rect 12002 2694 12012 2746
rect 12036 2694 12066 2746
rect 12066 2694 12078 2746
rect 12078 2694 12092 2746
rect 12116 2694 12130 2746
rect 12130 2694 12142 2746
rect 12142 2694 12172 2746
rect 12196 2694 12206 2746
rect 12206 2694 12252 2746
rect 11956 2692 12012 2694
rect 12036 2692 12092 2694
rect 12116 2692 12172 2694
rect 12196 2692 12252 2694
rect 14094 8336 14150 8392
rect 14094 5208 14150 5264
rect 14830 15000 14886 15056
rect 14830 13640 14886 13696
rect 14830 11212 14886 11248
rect 14830 11192 14832 11212
rect 14832 11192 14884 11212
rect 14884 11192 14886 11212
rect 14370 3440 14426 3496
rect 15106 10920 15162 10976
rect 15658 13504 15714 13560
rect 15382 11056 15438 11112
rect 15014 10240 15070 10296
rect 14830 5752 14886 5808
rect 15198 9696 15254 9752
rect 15106 8880 15162 8936
rect 15198 8472 15254 8528
rect 15106 6840 15162 6896
rect 15382 8200 15438 8256
rect 15382 4664 15438 4720
rect 15842 13368 15898 13424
rect 15658 11464 15714 11520
rect 15750 9696 15806 9752
rect 15658 7248 15714 7304
rect 15934 11056 15990 11112
rect 16118 12960 16174 13016
rect 16210 11056 16266 11112
rect 17616 17434 17672 17436
rect 17696 17434 17752 17436
rect 17776 17434 17832 17436
rect 17856 17434 17912 17436
rect 17616 17382 17662 17434
rect 17662 17382 17672 17434
rect 17696 17382 17726 17434
rect 17726 17382 17738 17434
rect 17738 17382 17752 17434
rect 17776 17382 17790 17434
rect 17790 17382 17802 17434
rect 17802 17382 17832 17434
rect 17856 17382 17866 17434
rect 17866 17382 17912 17434
rect 17616 17380 17672 17382
rect 17696 17380 17752 17382
rect 17776 17380 17832 17382
rect 17856 17380 17912 17382
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 17002 16890
rect 17002 16838 17012 16890
rect 17036 16838 17066 16890
rect 17066 16838 17078 16890
rect 17078 16838 17092 16890
rect 17116 16838 17130 16890
rect 17130 16838 17142 16890
rect 17142 16838 17172 16890
rect 17196 16838 17206 16890
rect 17206 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16394 11600 16450 11656
rect 16394 11056 16450 11112
rect 16486 10512 16542 10568
rect 16302 9560 16358 9616
rect 16118 6704 16174 6760
rect 16578 9968 16634 10024
rect 16946 15952 17002 16008
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 17002 15802
rect 17002 15750 17012 15802
rect 17036 15750 17066 15802
rect 17066 15750 17078 15802
rect 17078 15750 17092 15802
rect 17116 15750 17130 15802
rect 17130 15750 17142 15802
rect 17142 15750 17172 15802
rect 17196 15750 17206 15802
rect 17206 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16854 15544 16910 15600
rect 16854 15428 16910 15464
rect 16854 15408 16856 15428
rect 16856 15408 16908 15428
rect 16908 15408 16910 15428
rect 16762 14728 16818 14784
rect 16762 12824 16818 12880
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 17002 14714
rect 17002 14662 17012 14714
rect 17036 14662 17066 14714
rect 17066 14662 17078 14714
rect 17078 14662 17092 14714
rect 17116 14662 17130 14714
rect 17130 14662 17142 14714
rect 17142 14662 17172 14714
rect 17196 14662 17206 14714
rect 17206 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 17038 13912 17094 13968
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 17002 13626
rect 17002 13574 17012 13626
rect 17036 13574 17066 13626
rect 17066 13574 17078 13626
rect 17078 13574 17092 13626
rect 17116 13574 17130 13626
rect 17130 13574 17142 13626
rect 17142 13574 17172 13626
rect 17196 13574 17206 13626
rect 17206 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 17616 16346 17672 16348
rect 17696 16346 17752 16348
rect 17776 16346 17832 16348
rect 17856 16346 17912 16348
rect 17616 16294 17662 16346
rect 17662 16294 17672 16346
rect 17696 16294 17726 16346
rect 17726 16294 17738 16346
rect 17738 16294 17752 16346
rect 17776 16294 17790 16346
rect 17790 16294 17802 16346
rect 17802 16294 17832 16346
rect 17856 16294 17866 16346
rect 17866 16294 17912 16346
rect 17616 16292 17672 16294
rect 17696 16292 17752 16294
rect 17776 16292 17832 16294
rect 17856 16292 17912 16294
rect 17498 16088 17554 16144
rect 17616 15258 17672 15260
rect 17696 15258 17752 15260
rect 17776 15258 17832 15260
rect 17856 15258 17912 15260
rect 17616 15206 17662 15258
rect 17662 15206 17672 15258
rect 17696 15206 17726 15258
rect 17726 15206 17738 15258
rect 17738 15206 17752 15258
rect 17776 15206 17790 15258
rect 17790 15206 17802 15258
rect 17802 15206 17832 15258
rect 17856 15206 17866 15258
rect 17866 15206 17912 15258
rect 17616 15204 17672 15206
rect 17696 15204 17752 15206
rect 17776 15204 17832 15206
rect 17856 15204 17912 15206
rect 17616 14170 17672 14172
rect 17696 14170 17752 14172
rect 17776 14170 17832 14172
rect 17856 14170 17912 14172
rect 17616 14118 17662 14170
rect 17662 14118 17672 14170
rect 17696 14118 17726 14170
rect 17726 14118 17738 14170
rect 17738 14118 17752 14170
rect 17776 14118 17790 14170
rect 17790 14118 17802 14170
rect 17802 14118 17832 14170
rect 17856 14118 17866 14170
rect 17866 14118 17912 14170
rect 17616 14116 17672 14118
rect 17696 14116 17752 14118
rect 17776 14116 17832 14118
rect 17856 14116 17912 14118
rect 17616 13082 17672 13084
rect 17696 13082 17752 13084
rect 17776 13082 17832 13084
rect 17856 13082 17912 13084
rect 17616 13030 17662 13082
rect 17662 13030 17672 13082
rect 17696 13030 17726 13082
rect 17726 13030 17738 13082
rect 17738 13030 17752 13082
rect 17776 13030 17790 13082
rect 17790 13030 17802 13082
rect 17802 13030 17832 13082
rect 17856 13030 17866 13082
rect 17866 13030 17912 13082
rect 17616 13028 17672 13030
rect 17696 13028 17752 13030
rect 17776 13028 17832 13030
rect 17856 13028 17912 13030
rect 16854 12688 16910 12744
rect 17314 12688 17370 12744
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 17002 12538
rect 17002 12486 17012 12538
rect 17036 12486 17066 12538
rect 17066 12486 17078 12538
rect 17078 12486 17092 12538
rect 17116 12486 17130 12538
rect 17130 12486 17142 12538
rect 17142 12486 17172 12538
rect 17196 12486 17206 12538
rect 17206 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 17406 12280 17462 12336
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 17002 11450
rect 17002 11398 17012 11450
rect 17036 11398 17066 11450
rect 17066 11398 17078 11450
rect 17078 11398 17092 11450
rect 17116 11398 17130 11450
rect 17130 11398 17142 11450
rect 17142 11398 17172 11450
rect 17196 11398 17206 11450
rect 17206 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 17002 10362
rect 17002 10310 17012 10362
rect 17036 10310 17066 10362
rect 17066 10310 17078 10362
rect 17078 10310 17092 10362
rect 17116 10310 17130 10362
rect 17130 10310 17142 10362
rect 17142 10310 17172 10362
rect 17196 10310 17206 10362
rect 17206 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 17130 9460 17132 9480
rect 17132 9460 17184 9480
rect 17184 9460 17186 9480
rect 17130 9424 17186 9460
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 17002 9274
rect 17002 9222 17012 9274
rect 17036 9222 17066 9274
rect 17066 9222 17078 9274
rect 17078 9222 17092 9274
rect 17116 9222 17130 9274
rect 17130 9222 17142 9274
rect 17142 9222 17172 9274
rect 17196 9222 17206 9274
rect 17206 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 17002 8186
rect 17002 8134 17012 8186
rect 17036 8134 17066 8186
rect 17066 8134 17078 8186
rect 17078 8134 17092 8186
rect 17116 8134 17130 8186
rect 17130 8134 17142 8186
rect 17142 8134 17172 8186
rect 17196 8134 17206 8186
rect 17206 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 16762 5888 16818 5944
rect 15658 4564 15660 4584
rect 15660 4564 15712 4584
rect 15712 4564 15714 4584
rect 15658 4528 15714 4564
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 17002 7098
rect 17002 7046 17012 7098
rect 17036 7046 17066 7098
rect 17066 7046 17078 7098
rect 17078 7046 17092 7098
rect 17116 7046 17130 7098
rect 17130 7046 17142 7098
rect 17142 7046 17172 7098
rect 17196 7046 17206 7098
rect 17206 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 17002 6010
rect 17002 5958 17012 6010
rect 17036 5958 17066 6010
rect 17066 5958 17078 6010
rect 17078 5958 17092 6010
rect 17116 5958 17130 6010
rect 17130 5958 17142 6010
rect 17142 5958 17172 6010
rect 17196 5958 17206 6010
rect 17206 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 17002 4922
rect 17002 4870 17012 4922
rect 17036 4870 17066 4922
rect 17066 4870 17078 4922
rect 17078 4870 17092 4922
rect 17116 4870 17130 4922
rect 17130 4870 17142 4922
rect 17142 4870 17172 4922
rect 17196 4870 17206 4922
rect 17206 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 15750 2488 15806 2544
rect 16118 2372 16174 2408
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 17002 3834
rect 17002 3782 17012 3834
rect 17036 3782 17066 3834
rect 17066 3782 17078 3834
rect 17078 3782 17092 3834
rect 17116 3782 17130 3834
rect 17130 3782 17142 3834
rect 17142 3782 17172 3834
rect 17196 3782 17206 3834
rect 17206 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 17002 2746
rect 17002 2694 17012 2746
rect 17036 2694 17066 2746
rect 17066 2694 17078 2746
rect 17078 2694 17092 2746
rect 17116 2694 17130 2746
rect 17130 2694 17142 2746
rect 17142 2694 17172 2746
rect 17196 2694 17206 2746
rect 17206 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 17616 11994 17672 11996
rect 17696 11994 17752 11996
rect 17776 11994 17832 11996
rect 17856 11994 17912 11996
rect 17616 11942 17662 11994
rect 17662 11942 17672 11994
rect 17696 11942 17726 11994
rect 17726 11942 17738 11994
rect 17738 11942 17752 11994
rect 17776 11942 17790 11994
rect 17790 11942 17802 11994
rect 17802 11942 17832 11994
rect 17856 11942 17866 11994
rect 17866 11942 17912 11994
rect 17616 11940 17672 11942
rect 17696 11940 17752 11942
rect 17776 11940 17832 11942
rect 17856 11940 17912 11942
rect 17616 10906 17672 10908
rect 17696 10906 17752 10908
rect 17776 10906 17832 10908
rect 17856 10906 17912 10908
rect 17616 10854 17662 10906
rect 17662 10854 17672 10906
rect 17696 10854 17726 10906
rect 17726 10854 17738 10906
rect 17738 10854 17752 10906
rect 17776 10854 17790 10906
rect 17790 10854 17802 10906
rect 17802 10854 17832 10906
rect 17856 10854 17866 10906
rect 17866 10854 17912 10906
rect 17616 10852 17672 10854
rect 17696 10852 17752 10854
rect 17776 10852 17832 10854
rect 17856 10852 17912 10854
rect 17866 10124 17922 10160
rect 17866 10104 17868 10124
rect 17868 10104 17920 10124
rect 17920 10104 17922 10124
rect 17616 9818 17672 9820
rect 17696 9818 17752 9820
rect 17776 9818 17832 9820
rect 17856 9818 17912 9820
rect 17616 9766 17662 9818
rect 17662 9766 17672 9818
rect 17696 9766 17726 9818
rect 17726 9766 17738 9818
rect 17738 9766 17752 9818
rect 17776 9766 17790 9818
rect 17790 9766 17802 9818
rect 17802 9766 17832 9818
rect 17856 9766 17866 9818
rect 17866 9766 17912 9818
rect 17616 9764 17672 9766
rect 17696 9764 17752 9766
rect 17776 9764 17832 9766
rect 17856 9764 17912 9766
rect 17958 9016 18014 9072
rect 17616 8730 17672 8732
rect 17696 8730 17752 8732
rect 17776 8730 17832 8732
rect 17856 8730 17912 8732
rect 17616 8678 17662 8730
rect 17662 8678 17672 8730
rect 17696 8678 17726 8730
rect 17726 8678 17738 8730
rect 17738 8678 17752 8730
rect 17776 8678 17790 8730
rect 17790 8678 17802 8730
rect 17802 8678 17832 8730
rect 17856 8678 17866 8730
rect 17866 8678 17912 8730
rect 17616 8676 17672 8678
rect 17696 8676 17752 8678
rect 17776 8676 17832 8678
rect 17856 8676 17912 8678
rect 17682 7928 17738 7984
rect 17616 7642 17672 7644
rect 17696 7642 17752 7644
rect 17776 7642 17832 7644
rect 17856 7642 17912 7644
rect 17616 7590 17662 7642
rect 17662 7590 17672 7642
rect 17696 7590 17726 7642
rect 17726 7590 17738 7642
rect 17738 7590 17752 7642
rect 17776 7590 17790 7642
rect 17790 7590 17802 7642
rect 17802 7590 17832 7642
rect 17856 7590 17866 7642
rect 17866 7590 17912 7642
rect 17616 7588 17672 7590
rect 17696 7588 17752 7590
rect 17776 7588 17832 7590
rect 17856 7588 17912 7590
rect 17616 6554 17672 6556
rect 17696 6554 17752 6556
rect 17776 6554 17832 6556
rect 17856 6554 17912 6556
rect 17616 6502 17662 6554
rect 17662 6502 17672 6554
rect 17696 6502 17726 6554
rect 17726 6502 17738 6554
rect 17738 6502 17752 6554
rect 17776 6502 17790 6554
rect 17790 6502 17802 6554
rect 17802 6502 17832 6554
rect 17856 6502 17866 6554
rect 17866 6502 17912 6554
rect 17616 6500 17672 6502
rect 17696 6500 17752 6502
rect 17776 6500 17832 6502
rect 17856 6500 17912 6502
rect 17616 5466 17672 5468
rect 17696 5466 17752 5468
rect 17776 5466 17832 5468
rect 17856 5466 17912 5468
rect 17616 5414 17662 5466
rect 17662 5414 17672 5466
rect 17696 5414 17726 5466
rect 17726 5414 17738 5466
rect 17738 5414 17752 5466
rect 17776 5414 17790 5466
rect 17790 5414 17802 5466
rect 17802 5414 17832 5466
rect 17856 5414 17866 5466
rect 17866 5414 17912 5466
rect 17616 5412 17672 5414
rect 17696 5412 17752 5414
rect 17776 5412 17832 5414
rect 17856 5412 17912 5414
rect 17616 4378 17672 4380
rect 17696 4378 17752 4380
rect 17776 4378 17832 4380
rect 17856 4378 17912 4380
rect 17616 4326 17662 4378
rect 17662 4326 17672 4378
rect 17696 4326 17726 4378
rect 17726 4326 17738 4378
rect 17738 4326 17752 4378
rect 17776 4326 17790 4378
rect 17790 4326 17802 4378
rect 17802 4326 17832 4378
rect 17856 4326 17866 4378
rect 17866 4326 17912 4378
rect 17616 4324 17672 4326
rect 17696 4324 17752 4326
rect 17776 4324 17832 4326
rect 17856 4324 17912 4326
rect 17616 3290 17672 3292
rect 17696 3290 17752 3292
rect 17776 3290 17832 3292
rect 17856 3290 17912 3292
rect 17616 3238 17662 3290
rect 17662 3238 17672 3290
rect 17696 3238 17726 3290
rect 17726 3238 17738 3290
rect 17738 3238 17752 3290
rect 17776 3238 17790 3290
rect 17790 3238 17802 3290
rect 17802 3238 17832 3290
rect 17856 3238 17866 3290
rect 17866 3238 17912 3290
rect 17616 3236 17672 3238
rect 17696 3236 17752 3238
rect 17776 3236 17832 3238
rect 17856 3236 17912 3238
rect 16118 2352 16120 2372
rect 16120 2352 16172 2372
rect 16172 2352 16174 2372
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1858 1672 1914 1728
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 18418 13640 18474 13696
rect 18418 11192 18474 11248
rect 18418 8780 18420 8800
rect 18420 8780 18472 8800
rect 18472 8780 18474 8800
rect 18418 8744 18474 8780
rect 18234 6296 18290 6352
rect 18418 6296 18474 6352
rect 18418 3884 18420 3904
rect 18420 3884 18472 3904
rect 18472 3884 18474 3904
rect 18418 3848 18474 3884
rect 17616 2202 17672 2204
rect 17696 2202 17752 2204
rect 17776 2202 17832 2204
rect 17856 2202 17912 2204
rect 17616 2150 17662 2202
rect 17662 2150 17672 2202
rect 17696 2150 17726 2202
rect 17726 2150 17738 2202
rect 17738 2150 17752 2202
rect 17776 2150 17790 2202
rect 17790 2150 17802 2202
rect 17802 2150 17832 2202
rect 17856 2150 17866 2202
rect 17866 2150 17912 2202
rect 17616 2148 17672 2150
rect 17696 2148 17752 2150
rect 17776 2148 17832 2150
rect 17856 2148 17912 2150
rect 18418 1400 18474 1456
<< metal3 >>
rect 17861 18594 17927 18597
rect 19200 18594 20000 18624
rect 17861 18592 20000 18594
rect 17861 18536 17866 18592
rect 17922 18536 20000 18592
rect 17861 18534 20000 18536
rect 17861 18531 17927 18534
rect 19200 18504 20000 18534
rect 0 18050 800 18080
rect 1853 18050 1919 18053
rect 0 18048 1919 18050
rect 0 17992 1858 18048
rect 1914 17992 1919 18048
rect 0 17990 1919 17992
rect 0 17960 800 17990
rect 1853 17987 1919 17990
rect 2606 17440 2922 17441
rect 2606 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2922 17440
rect 2606 17375 2922 17376
rect 7606 17440 7922 17441
rect 7606 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7922 17440
rect 7606 17375 7922 17376
rect 12606 17440 12922 17441
rect 12606 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12922 17440
rect 12606 17375 12922 17376
rect 17606 17440 17922 17441
rect 17606 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17922 17440
rect 17606 17375 17922 17376
rect 841 17098 907 17101
rect 798 17096 907 17098
rect 798 17040 846 17096
rect 902 17040 907 17096
rect 798 17035 907 17040
rect 5942 17036 5948 17100
rect 6012 17098 6018 17100
rect 14089 17098 14155 17101
rect 6012 17096 14155 17098
rect 6012 17040 14094 17096
rect 14150 17040 14155 17096
rect 6012 17038 14155 17040
rect 6012 17036 6018 17038
rect 14089 17035 14155 17038
rect 798 16992 858 17035
rect 0 16902 858 16992
rect 0 16872 800 16902
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 6946 16896 7262 16897
rect 6946 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7262 16896
rect 6946 16831 7262 16832
rect 11946 16896 12262 16897
rect 11946 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12262 16896
rect 11946 16831 12262 16832
rect 16946 16896 17262 16897
rect 16946 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17262 16896
rect 16946 16831 17262 16832
rect 11094 16628 11100 16692
rect 11164 16690 11170 16692
rect 15193 16690 15259 16693
rect 11164 16688 15259 16690
rect 11164 16632 15198 16688
rect 15254 16632 15259 16688
rect 11164 16630 15259 16632
rect 11164 16628 11170 16630
rect 15193 16627 15259 16630
rect 6913 16554 6979 16557
rect 10317 16554 10383 16557
rect 14181 16554 14247 16557
rect 6913 16552 10383 16554
rect 6913 16496 6918 16552
rect 6974 16496 10322 16552
rect 10378 16496 10383 16552
rect 6913 16494 10383 16496
rect 6913 16491 6979 16494
rect 10317 16491 10383 16494
rect 12390 16552 14247 16554
rect 12390 16496 14186 16552
rect 14242 16496 14247 16552
rect 12390 16494 14247 16496
rect 4705 16418 4771 16421
rect 7465 16418 7531 16421
rect 4705 16416 7531 16418
rect 4705 16360 4710 16416
rect 4766 16360 7470 16416
rect 7526 16360 7531 16416
rect 4705 16358 7531 16360
rect 4705 16355 4771 16358
rect 7465 16355 7531 16358
rect 8017 16418 8083 16421
rect 12390 16418 12450 16494
rect 14181 16491 14247 16494
rect 8017 16416 12450 16418
rect 8017 16360 8022 16416
rect 8078 16360 12450 16416
rect 8017 16358 12450 16360
rect 13261 16418 13327 16421
rect 14406 16418 14412 16420
rect 13261 16416 14412 16418
rect 13261 16360 13266 16416
rect 13322 16360 14412 16416
rect 13261 16358 14412 16360
rect 8017 16355 8083 16358
rect 13261 16355 13327 16358
rect 14406 16356 14412 16358
rect 14476 16356 14482 16420
rect 2606 16352 2922 16353
rect 2606 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2922 16352
rect 2606 16287 2922 16288
rect 7606 16352 7922 16353
rect 7606 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7922 16352
rect 7606 16287 7922 16288
rect 12606 16352 12922 16353
rect 12606 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12922 16352
rect 12606 16287 12922 16288
rect 17606 16352 17922 16353
rect 17606 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17922 16352
rect 17606 16287 17922 16288
rect 9397 16282 9463 16285
rect 11973 16282 12039 16285
rect 9397 16280 12039 16282
rect 9397 16224 9402 16280
rect 9458 16224 11978 16280
rect 12034 16224 12039 16280
rect 9397 16222 12039 16224
rect 9397 16219 9463 16222
rect 11973 16219 12039 16222
rect 12249 16146 12315 16149
rect 2730 16144 12315 16146
rect 2730 16088 12254 16144
rect 12310 16088 12315 16144
rect 2730 16086 12315 16088
rect 1485 16010 1551 16013
rect 2730 16010 2790 16086
rect 12249 16083 12315 16086
rect 17493 16146 17559 16149
rect 19200 16146 20000 16176
rect 17493 16144 20000 16146
rect 17493 16088 17498 16144
rect 17554 16088 20000 16144
rect 17493 16086 20000 16088
rect 17493 16083 17559 16086
rect 19200 16056 20000 16086
rect 1485 16008 2790 16010
rect 1485 15952 1490 16008
rect 1546 15952 2790 16008
rect 1485 15950 2790 15952
rect 3049 16010 3115 16013
rect 4654 16010 4660 16012
rect 3049 16008 4660 16010
rect 3049 15952 3054 16008
rect 3110 15952 4660 16008
rect 3049 15950 4660 15952
rect 1485 15947 1551 15950
rect 3049 15947 3115 15950
rect 4654 15948 4660 15950
rect 4724 15948 4730 16012
rect 4797 16010 4863 16013
rect 5349 16010 5415 16013
rect 13629 16010 13695 16013
rect 16941 16010 17007 16013
rect 4797 16008 12450 16010
rect 4797 15952 4802 16008
rect 4858 15952 5354 16008
rect 5410 15952 12450 16008
rect 4797 15950 12450 15952
rect 4797 15947 4863 15950
rect 5349 15947 5415 15950
rect 0 15874 800 15904
rect 1025 15874 1091 15877
rect 0 15872 1091 15874
rect 0 15816 1030 15872
rect 1086 15816 1091 15872
rect 0 15814 1091 15816
rect 0 15784 800 15814
rect 1025 15811 1091 15814
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 6946 15808 7262 15809
rect 6946 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7262 15808
rect 6946 15743 7262 15744
rect 11946 15808 12262 15809
rect 11946 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12262 15808
rect 11946 15743 12262 15744
rect 10041 15738 10107 15741
rect 7422 15736 10107 15738
rect 7422 15680 10046 15736
rect 10102 15680 10107 15736
rect 7422 15678 10107 15680
rect 4337 15602 4403 15605
rect 7422 15602 7482 15678
rect 10041 15675 10107 15678
rect 4337 15600 7482 15602
rect 4337 15544 4342 15600
rect 4398 15544 7482 15600
rect 4337 15542 7482 15544
rect 9029 15602 9095 15605
rect 9254 15602 9260 15604
rect 9029 15600 9260 15602
rect 9029 15544 9034 15600
rect 9090 15544 9260 15600
rect 9029 15542 9260 15544
rect 4337 15539 4403 15542
rect 9029 15539 9095 15542
rect 9254 15540 9260 15542
rect 9324 15540 9330 15604
rect 12390 15602 12450 15950
rect 13629 16008 17007 16010
rect 13629 15952 13634 16008
rect 13690 15952 16946 16008
rect 17002 15952 17007 16008
rect 13629 15950 17007 15952
rect 13629 15947 13695 15950
rect 16941 15947 17007 15950
rect 16946 15808 17262 15809
rect 16946 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17262 15808
rect 16946 15743 17262 15744
rect 13537 15602 13603 15605
rect 12390 15600 13603 15602
rect 12390 15544 13542 15600
rect 13598 15544 13603 15600
rect 12390 15542 13603 15544
rect 13537 15539 13603 15542
rect 16614 15540 16620 15604
rect 16684 15602 16690 15604
rect 16849 15602 16915 15605
rect 16684 15600 16915 15602
rect 16684 15544 16854 15600
rect 16910 15544 16915 15600
rect 16684 15542 16915 15544
rect 16684 15540 16690 15542
rect 16849 15539 16915 15542
rect 6494 15404 6500 15468
rect 6564 15466 6570 15468
rect 9121 15466 9187 15469
rect 6564 15464 9187 15466
rect 6564 15408 9126 15464
rect 9182 15408 9187 15464
rect 6564 15406 9187 15408
rect 6564 15404 6570 15406
rect 9121 15403 9187 15406
rect 9765 15466 9831 15469
rect 10685 15466 10751 15469
rect 9765 15464 10751 15466
rect 9765 15408 9770 15464
rect 9826 15408 10690 15464
rect 10746 15408 10751 15464
rect 9765 15406 10751 15408
rect 9765 15403 9831 15406
rect 10685 15403 10751 15406
rect 11421 15466 11487 15469
rect 16849 15466 16915 15469
rect 11421 15464 16915 15466
rect 11421 15408 11426 15464
rect 11482 15408 16854 15464
rect 16910 15408 16915 15464
rect 11421 15406 16915 15408
rect 11421 15403 11487 15406
rect 16849 15403 16915 15406
rect 6637 15332 6703 15333
rect 9397 15332 9463 15333
rect 10409 15332 10475 15333
rect 6637 15328 6684 15332
rect 6748 15330 6754 15332
rect 6637 15272 6642 15328
rect 6637 15268 6684 15272
rect 6748 15270 6794 15330
rect 9397 15328 9444 15332
rect 9508 15330 9514 15332
rect 10358 15330 10364 15332
rect 9397 15272 9402 15328
rect 6748 15268 6754 15270
rect 9397 15268 9444 15272
rect 9508 15270 9554 15330
rect 10318 15270 10364 15330
rect 10428 15328 10475 15332
rect 10470 15272 10475 15328
rect 9508 15268 9514 15270
rect 10358 15268 10364 15270
rect 10428 15268 10475 15272
rect 6637 15267 6703 15268
rect 9397 15267 9463 15268
rect 10409 15267 10475 15268
rect 10593 15330 10659 15333
rect 10961 15332 11027 15333
rect 10726 15330 10732 15332
rect 10593 15328 10732 15330
rect 10593 15272 10598 15328
rect 10654 15272 10732 15328
rect 10593 15270 10732 15272
rect 10593 15267 10659 15270
rect 10726 15268 10732 15270
rect 10796 15268 10802 15332
rect 10910 15330 10916 15332
rect 10870 15270 10916 15330
rect 10980 15328 11027 15332
rect 11022 15272 11027 15328
rect 10910 15268 10916 15270
rect 10980 15268 11027 15272
rect 10961 15267 11027 15268
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 7606 15264 7922 15265
rect 7606 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7922 15264
rect 7606 15199 7922 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 12606 15199 12922 15200
rect 17606 15264 17922 15265
rect 17606 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17922 15264
rect 17606 15199 17922 15200
rect 9673 15194 9739 15197
rect 10317 15194 10383 15197
rect 10961 15194 11027 15197
rect 9673 15192 11027 15194
rect 9673 15136 9678 15192
rect 9734 15136 10322 15192
rect 10378 15136 10966 15192
rect 11022 15136 11027 15192
rect 9673 15134 11027 15136
rect 9673 15131 9739 15134
rect 10317 15131 10383 15134
rect 10961 15131 11027 15134
rect 3969 15058 4035 15061
rect 10133 15058 10199 15061
rect 14825 15058 14891 15061
rect 3969 15056 14891 15058
rect 3969 15000 3974 15056
rect 4030 15000 10138 15056
rect 10194 15000 14830 15056
rect 14886 15000 14891 15056
rect 3969 14998 14891 15000
rect 3969 14995 4035 14998
rect 10133 14995 10199 14998
rect 14825 14995 14891 14998
rect 841 14922 907 14925
rect 798 14920 907 14922
rect 798 14864 846 14920
rect 902 14864 907 14920
rect 798 14859 907 14864
rect 9765 14922 9831 14925
rect 14365 14922 14431 14925
rect 9765 14920 14431 14922
rect 9765 14864 9770 14920
rect 9826 14864 14370 14920
rect 14426 14864 14431 14920
rect 9765 14862 14431 14864
rect 9765 14859 9831 14862
rect 14365 14859 14431 14862
rect 798 14816 858 14859
rect 0 14726 858 14816
rect 9673 14786 9739 14789
rect 10593 14788 10659 14789
rect 9806 14786 9812 14788
rect 9673 14784 9812 14786
rect 9673 14728 9678 14784
rect 9734 14728 9812 14784
rect 9673 14726 9812 14728
rect 0 14696 800 14726
rect 9673 14723 9739 14726
rect 9806 14724 9812 14726
rect 9876 14724 9882 14788
rect 10542 14724 10548 14788
rect 10612 14786 10659 14788
rect 12341 14786 12407 14789
rect 16757 14786 16823 14789
rect 10612 14784 10704 14786
rect 10654 14728 10704 14784
rect 10612 14726 10704 14728
rect 12341 14784 16823 14786
rect 12341 14728 12346 14784
rect 12402 14728 16762 14784
rect 16818 14728 16823 14784
rect 12341 14726 16823 14728
rect 10612 14724 10659 14726
rect 10593 14723 10659 14724
rect 12341 14723 12407 14726
rect 16757 14723 16823 14726
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 6946 14720 7262 14721
rect 6946 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7262 14720
rect 6946 14655 7262 14656
rect 11946 14720 12262 14721
rect 11946 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12262 14720
rect 11946 14655 12262 14656
rect 16946 14720 17262 14721
rect 16946 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17262 14720
rect 16946 14655 17262 14656
rect 9673 14650 9739 14653
rect 10501 14650 10567 14653
rect 9673 14648 10567 14650
rect 9673 14592 9678 14648
rect 9734 14592 10506 14648
rect 10562 14592 10567 14648
rect 9673 14590 10567 14592
rect 9673 14587 9739 14590
rect 10501 14587 10567 14590
rect 12525 14650 12591 14653
rect 14273 14650 14339 14653
rect 12525 14648 14339 14650
rect 12525 14592 12530 14648
rect 12586 14592 14278 14648
rect 14334 14592 14339 14648
rect 12525 14590 14339 14592
rect 12525 14587 12591 14590
rect 14273 14587 14339 14590
rect 6821 14514 6887 14517
rect 9765 14514 9831 14517
rect 6821 14512 9831 14514
rect 6821 14456 6826 14512
rect 6882 14456 9770 14512
rect 9826 14456 9831 14512
rect 6821 14454 9831 14456
rect 6821 14451 6887 14454
rect 9765 14451 9831 14454
rect 9990 14452 9996 14516
rect 10060 14514 10066 14516
rect 10593 14514 10659 14517
rect 14549 14514 14615 14517
rect 10060 14512 14615 14514
rect 10060 14456 10598 14512
rect 10654 14456 14554 14512
rect 14610 14456 14615 14512
rect 10060 14454 14615 14456
rect 10060 14452 10066 14454
rect 10593 14451 10659 14454
rect 14549 14451 14615 14454
rect 3918 14316 3924 14380
rect 3988 14378 3994 14380
rect 9581 14378 9647 14381
rect 15326 14378 15332 14380
rect 3988 14318 8218 14378
rect 3988 14316 3994 14318
rect 8158 14242 8218 14318
rect 9581 14376 15332 14378
rect 9581 14320 9586 14376
rect 9642 14320 15332 14376
rect 9581 14318 15332 14320
rect 9581 14315 9647 14318
rect 15326 14316 15332 14318
rect 15396 14316 15402 14380
rect 11421 14242 11487 14245
rect 8158 14240 11487 14242
rect 8158 14184 11426 14240
rect 11482 14184 11487 14240
rect 8158 14182 11487 14184
rect 11421 14179 11487 14182
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 7606 14176 7922 14177
rect 7606 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7922 14176
rect 7606 14111 7922 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 12606 14111 12922 14112
rect 17606 14176 17922 14177
rect 17606 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17922 14176
rect 17606 14111 17922 14112
rect 8150 13908 8156 13972
rect 8220 13970 8226 13972
rect 10133 13970 10199 13973
rect 8220 13968 10199 13970
rect 8220 13912 10138 13968
rect 10194 13912 10199 13968
rect 8220 13910 10199 13912
rect 8220 13908 8226 13910
rect 10133 13907 10199 13910
rect 10317 13970 10383 13973
rect 17033 13970 17099 13973
rect 10317 13968 17099 13970
rect 10317 13912 10322 13968
rect 10378 13912 17038 13968
rect 17094 13912 17099 13968
rect 10317 13910 17099 13912
rect 10317 13907 10383 13910
rect 17033 13907 17099 13910
rect 3509 13834 3575 13837
rect 6126 13834 6132 13836
rect 3509 13832 6132 13834
rect 3509 13776 3514 13832
rect 3570 13776 6132 13832
rect 3509 13774 6132 13776
rect 3509 13771 3575 13774
rect 6126 13772 6132 13774
rect 6196 13772 6202 13836
rect 8661 13834 8727 13837
rect 9121 13834 9187 13837
rect 8661 13832 9187 13834
rect 8661 13776 8666 13832
rect 8722 13776 9126 13832
rect 9182 13776 9187 13832
rect 8661 13774 9187 13776
rect 8661 13771 8727 13774
rect 9121 13771 9187 13774
rect 11654 13774 12450 13834
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 6946 13632 7262 13633
rect 6946 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7262 13632
rect 6946 13567 7262 13568
rect 9070 13500 9076 13564
rect 9140 13562 9146 13564
rect 11654 13562 11714 13774
rect 12390 13698 12450 13774
rect 13486 13772 13492 13836
rect 13556 13834 13562 13836
rect 13629 13834 13695 13837
rect 13556 13832 13695 13834
rect 13556 13776 13634 13832
rect 13690 13776 13695 13832
rect 13556 13774 13695 13776
rect 13556 13772 13562 13774
rect 13629 13771 13695 13774
rect 13813 13834 13879 13837
rect 14958 13834 14964 13836
rect 13813 13832 14964 13834
rect 13813 13776 13818 13832
rect 13874 13776 14964 13832
rect 13813 13774 14964 13776
rect 13813 13771 13879 13774
rect 14958 13772 14964 13774
rect 15028 13772 15034 13836
rect 12985 13698 13051 13701
rect 12390 13696 13051 13698
rect 12390 13640 12990 13696
rect 13046 13640 13051 13696
rect 12390 13638 13051 13640
rect 12985 13635 13051 13638
rect 13445 13698 13511 13701
rect 14825 13698 14891 13701
rect 13445 13696 14891 13698
rect 13445 13640 13450 13696
rect 13506 13640 14830 13696
rect 14886 13640 14891 13696
rect 13445 13638 14891 13640
rect 13445 13635 13511 13638
rect 14825 13635 14891 13638
rect 18413 13698 18479 13701
rect 19200 13698 20000 13728
rect 18413 13696 20000 13698
rect 18413 13640 18418 13696
rect 18474 13640 20000 13696
rect 18413 13638 20000 13640
rect 18413 13635 18479 13638
rect 11946 13632 12262 13633
rect 11946 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12262 13632
rect 11946 13567 12262 13568
rect 16946 13632 17262 13633
rect 16946 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17262 13632
rect 19200 13608 20000 13638
rect 16946 13567 17262 13568
rect 15653 13562 15719 13565
rect 15878 13562 15884 13564
rect 9140 13502 11714 13562
rect 12390 13560 15884 13562
rect 12390 13504 15658 13560
rect 15714 13504 15884 13560
rect 12390 13502 15884 13504
rect 9140 13500 9146 13502
rect 4889 13426 4955 13429
rect 8293 13426 8359 13429
rect 12390 13426 12450 13502
rect 15653 13499 15719 13502
rect 15878 13500 15884 13502
rect 15948 13500 15954 13564
rect 4889 13424 7804 13426
rect 4889 13368 4894 13424
rect 4950 13368 7804 13424
rect 4889 13366 7804 13368
rect 4889 13363 4955 13366
rect 7414 13228 7420 13292
rect 7484 13290 7490 13292
rect 7557 13290 7623 13293
rect 7484 13288 7623 13290
rect 7484 13232 7562 13288
rect 7618 13232 7623 13288
rect 7484 13230 7623 13232
rect 7744 13290 7804 13366
rect 8293 13424 12450 13426
rect 8293 13368 8298 13424
rect 8354 13368 12450 13424
rect 8293 13366 12450 13368
rect 12709 13426 12775 13429
rect 13670 13426 13676 13428
rect 12709 13424 13676 13426
rect 12709 13368 12714 13424
rect 12770 13368 13676 13424
rect 12709 13366 13676 13368
rect 8293 13363 8359 13366
rect 12709 13363 12775 13366
rect 13670 13364 13676 13366
rect 13740 13426 13746 13428
rect 15837 13426 15903 13429
rect 13740 13424 15903 13426
rect 13740 13368 15842 13424
rect 15898 13368 15903 13424
rect 13740 13366 15903 13368
rect 13740 13364 13746 13366
rect 15837 13363 15903 13366
rect 9581 13290 9647 13293
rect 14549 13290 14615 13293
rect 7744 13288 9647 13290
rect 7744 13232 9586 13288
rect 9642 13232 9647 13288
rect 7744 13230 9647 13232
rect 7484 13228 7490 13230
rect 7557 13227 7623 13230
rect 9581 13227 9647 13230
rect 12390 13288 14615 13290
rect 12390 13232 14554 13288
rect 14610 13232 14615 13288
rect 12390 13230 14615 13232
rect 9254 13092 9260 13156
rect 9324 13154 9330 13156
rect 12390 13154 12450 13230
rect 14549 13227 14615 13230
rect 9324 13094 12450 13154
rect 9324 13092 9330 13094
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 7606 13088 7922 13089
rect 7606 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7922 13088
rect 7606 13023 7922 13024
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 12606 13023 12922 13024
rect 17606 13088 17922 13089
rect 17606 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17922 13088
rect 17606 13023 17922 13024
rect 13077 13018 13143 13021
rect 16113 13018 16179 13021
rect 13077 13016 16179 13018
rect 13077 12960 13082 13016
rect 13138 12960 16118 13016
rect 16174 12960 16179 13016
rect 13077 12958 16179 12960
rect 13077 12955 13143 12958
rect 16113 12955 16179 12958
rect 4429 12882 4495 12885
rect 8661 12882 8727 12885
rect 4429 12880 8727 12882
rect 4429 12824 4434 12880
rect 4490 12824 8666 12880
rect 8722 12824 8727 12880
rect 4429 12822 8727 12824
rect 4429 12819 4495 12822
rect 8661 12819 8727 12822
rect 9857 12882 9923 12885
rect 13997 12882 14063 12885
rect 16757 12882 16823 12885
rect 9857 12880 14063 12882
rect 9857 12824 9862 12880
rect 9918 12824 14002 12880
rect 14058 12824 14063 12880
rect 9857 12822 14063 12824
rect 9857 12819 9923 12822
rect 13997 12819 14063 12822
rect 16622 12880 16823 12882
rect 16622 12824 16762 12880
rect 16818 12824 16823 12880
rect 16622 12822 16823 12824
rect 841 12746 907 12749
rect 798 12744 907 12746
rect 798 12688 846 12744
rect 902 12688 907 12744
rect 798 12683 907 12688
rect 5390 12684 5396 12748
rect 5460 12746 5466 12748
rect 7005 12746 7071 12749
rect 5460 12744 7071 12746
rect 5460 12688 7010 12744
rect 7066 12688 7071 12744
rect 5460 12686 7071 12688
rect 5460 12684 5466 12686
rect 7005 12683 7071 12686
rect 7189 12746 7255 12749
rect 8845 12746 8911 12749
rect 7189 12744 8911 12746
rect 7189 12688 7194 12744
rect 7250 12688 8850 12744
rect 8906 12688 8911 12744
rect 7189 12686 8911 12688
rect 7189 12683 7255 12686
rect 8845 12683 8911 12686
rect 9673 12746 9739 12749
rect 16622 12746 16682 12822
rect 16757 12819 16823 12822
rect 16849 12748 16915 12749
rect 9673 12744 16682 12746
rect 9673 12688 9678 12744
rect 9734 12688 16682 12744
rect 9673 12686 16682 12688
rect 9673 12683 9739 12686
rect 16798 12684 16804 12748
rect 16868 12746 16915 12748
rect 17309 12748 17375 12749
rect 16868 12744 16960 12746
rect 16910 12688 16960 12744
rect 16868 12686 16960 12688
rect 17309 12744 17356 12748
rect 17420 12746 17426 12748
rect 17309 12688 17314 12744
rect 16868 12684 16915 12686
rect 16849 12683 16915 12684
rect 17309 12684 17356 12688
rect 17420 12686 17466 12746
rect 17420 12684 17426 12686
rect 17309 12683 17375 12684
rect 798 12640 858 12683
rect 0 12550 858 12640
rect 7741 12610 7807 12613
rect 8385 12610 8451 12613
rect 7741 12608 8451 12610
rect 7741 12552 7746 12608
rect 7802 12552 8390 12608
rect 8446 12552 8451 12608
rect 7741 12550 8451 12552
rect 0 12520 800 12550
rect 7741 12547 7807 12550
rect 8385 12547 8451 12550
rect 11053 12610 11119 12613
rect 11237 12610 11303 12613
rect 11053 12608 11303 12610
rect 11053 12552 11058 12608
rect 11114 12552 11242 12608
rect 11298 12552 11303 12608
rect 11053 12550 11303 12552
rect 11053 12547 11119 12550
rect 11237 12547 11303 12550
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 6946 12544 7262 12545
rect 6946 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7262 12544
rect 6946 12479 7262 12480
rect 11946 12544 12262 12545
rect 11946 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12262 12544
rect 11946 12479 12262 12480
rect 16946 12544 17262 12545
rect 16946 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17262 12544
rect 16946 12479 17262 12480
rect 9489 12474 9555 12477
rect 12617 12474 12683 12477
rect 13445 12474 13511 12477
rect 7606 12472 11162 12474
rect 7606 12416 9494 12472
rect 9550 12416 11162 12472
rect 7606 12414 11162 12416
rect 7189 12202 7255 12205
rect 7606 12202 7666 12414
rect 9489 12411 9555 12414
rect 7741 12338 7807 12341
rect 8150 12338 8156 12340
rect 7741 12336 8156 12338
rect 7741 12280 7746 12336
rect 7802 12280 8156 12336
rect 7741 12278 8156 12280
rect 7741 12275 7807 12278
rect 8150 12276 8156 12278
rect 8220 12276 8226 12340
rect 8385 12338 8451 12341
rect 9673 12338 9739 12341
rect 8385 12336 9739 12338
rect 8385 12280 8390 12336
rect 8446 12280 9678 12336
rect 9734 12280 9739 12336
rect 8385 12278 9739 12280
rect 11102 12338 11162 12414
rect 12617 12472 13511 12474
rect 12617 12416 12622 12472
rect 12678 12416 13450 12472
rect 13506 12416 13511 12472
rect 12617 12414 13511 12416
rect 12617 12411 12683 12414
rect 13445 12411 13511 12414
rect 11697 12338 11763 12341
rect 11973 12338 12039 12341
rect 11102 12336 12039 12338
rect 11102 12280 11702 12336
rect 11758 12280 11978 12336
rect 12034 12280 12039 12336
rect 11102 12278 12039 12280
rect 8385 12275 8451 12278
rect 9673 12275 9739 12278
rect 11697 12275 11763 12278
rect 11973 12275 12039 12278
rect 12985 12338 13051 12341
rect 13261 12338 13327 12341
rect 17401 12340 17467 12341
rect 17350 12338 17356 12340
rect 12985 12336 13327 12338
rect 12985 12280 12990 12336
rect 13046 12280 13266 12336
rect 13322 12280 13327 12336
rect 12985 12278 13327 12280
rect 17310 12278 17356 12338
rect 17420 12336 17467 12340
rect 17462 12280 17467 12336
rect 12985 12275 13051 12278
rect 13261 12275 13327 12278
rect 17350 12276 17356 12278
rect 17420 12276 17467 12280
rect 17401 12275 17467 12276
rect 7189 12200 7666 12202
rect 7189 12144 7194 12200
rect 7250 12144 7666 12200
rect 7189 12142 7666 12144
rect 8293 12202 8359 12205
rect 8293 12200 13186 12202
rect 8293 12144 8298 12200
rect 8354 12144 13186 12200
rect 8293 12142 13186 12144
rect 7189 12139 7255 12142
rect 8293 12139 8359 12142
rect 13126 12066 13186 12142
rect 13445 12066 13511 12069
rect 13126 12064 13511 12066
rect 13126 12008 13450 12064
rect 13506 12008 13511 12064
rect 13126 12006 13511 12008
rect 13445 12003 13511 12006
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 7606 12000 7922 12001
rect 7606 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7922 12000
rect 7606 11935 7922 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 12606 11935 12922 11936
rect 17606 12000 17922 12001
rect 17606 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17922 12000
rect 17606 11935 17922 11936
rect 10358 11930 10364 11932
rect 9262 11870 10364 11930
rect 7281 11794 7347 11797
rect 9262 11794 9322 11870
rect 10358 11868 10364 11870
rect 10428 11930 10434 11932
rect 10501 11930 10567 11933
rect 10428 11928 10567 11930
rect 10428 11872 10506 11928
rect 10562 11872 10567 11928
rect 10428 11870 10567 11872
rect 10428 11868 10434 11870
rect 10501 11867 10567 11870
rect 11646 11868 11652 11932
rect 11716 11930 11722 11932
rect 11881 11930 11947 11933
rect 11716 11928 11947 11930
rect 11716 11872 11886 11928
rect 11942 11872 11947 11928
rect 11716 11870 11947 11872
rect 11716 11868 11722 11870
rect 11881 11867 11947 11870
rect 7281 11792 9322 11794
rect 7281 11736 7286 11792
rect 7342 11736 9322 11792
rect 7281 11734 9322 11736
rect 9489 11794 9555 11797
rect 9489 11792 13554 11794
rect 9489 11736 9494 11792
rect 9550 11736 13554 11792
rect 9489 11734 13554 11736
rect 7281 11731 7347 11734
rect 9489 11731 9555 11734
rect 841 11658 907 11661
rect 798 11656 907 11658
rect 798 11600 846 11656
rect 902 11600 907 11656
rect 798 11595 907 11600
rect 3969 11658 4035 11661
rect 7833 11658 7899 11661
rect 3969 11656 7899 11658
rect 3969 11600 3974 11656
rect 4030 11600 7838 11656
rect 7894 11600 7899 11656
rect 3969 11598 7899 11600
rect 3969 11595 4035 11598
rect 7833 11595 7899 11598
rect 8017 11658 8083 11661
rect 12985 11658 13051 11661
rect 8017 11656 13051 11658
rect 8017 11600 8022 11656
rect 8078 11600 12990 11656
rect 13046 11600 13051 11656
rect 8017 11598 13051 11600
rect 13494 11658 13554 11734
rect 16389 11658 16455 11661
rect 13494 11656 16455 11658
rect 13494 11600 16394 11656
rect 16450 11600 16455 11656
rect 13494 11598 16455 11600
rect 8017 11595 8083 11598
rect 12985 11595 13051 11598
rect 16389 11595 16455 11598
rect 798 11552 858 11595
rect 0 11462 858 11552
rect 12709 11522 12775 11525
rect 15653 11522 15719 11525
rect 12709 11520 15719 11522
rect 12709 11464 12714 11520
rect 12770 11464 15658 11520
rect 15714 11464 15719 11520
rect 12709 11462 15719 11464
rect 0 11432 800 11462
rect 12709 11459 12775 11462
rect 15653 11459 15719 11462
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 11946 11456 12262 11457
rect 11946 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12262 11456
rect 11946 11391 12262 11392
rect 16946 11456 17262 11457
rect 16946 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17262 11456
rect 16946 11391 17262 11392
rect 5349 11386 5415 11389
rect 6729 11386 6795 11389
rect 5349 11384 6795 11386
rect 5349 11328 5354 11384
rect 5410 11328 6734 11384
rect 6790 11328 6795 11384
rect 5349 11326 6795 11328
rect 5349 11323 5415 11326
rect 6729 11323 6795 11326
rect 11094 11324 11100 11388
rect 11164 11386 11170 11388
rect 11513 11386 11579 11389
rect 11164 11384 11579 11386
rect 11164 11328 11518 11384
rect 11574 11328 11579 11384
rect 11164 11326 11579 11328
rect 11164 11324 11170 11326
rect 11513 11323 11579 11326
rect 14181 11386 14247 11389
rect 14181 11384 15578 11386
rect 14181 11328 14186 11384
rect 14242 11328 15578 11384
rect 14181 11326 15578 11328
rect 14181 11323 14247 11326
rect 1301 11250 1367 11253
rect 14825 11250 14891 11253
rect 1301 11248 14891 11250
rect 1301 11192 1306 11248
rect 1362 11192 14830 11248
rect 14886 11192 14891 11248
rect 1301 11190 14891 11192
rect 1301 11187 1367 11190
rect 14825 11187 14891 11190
rect 6453 11114 6519 11117
rect 15377 11114 15443 11117
rect 6453 11112 15443 11114
rect 6453 11056 6458 11112
rect 6514 11056 15382 11112
rect 15438 11056 15443 11112
rect 6453 11054 15443 11056
rect 15518 11114 15578 11326
rect 18413 11250 18479 11253
rect 19200 11250 20000 11280
rect 18413 11248 20000 11250
rect 18413 11192 18418 11248
rect 18474 11192 20000 11248
rect 18413 11190 20000 11192
rect 18413 11187 18479 11190
rect 19200 11160 20000 11190
rect 15929 11114 15995 11117
rect 15518 11112 15995 11114
rect 15518 11056 15934 11112
rect 15990 11056 15995 11112
rect 15518 11054 15995 11056
rect 6453 11051 6519 11054
rect 15377 11051 15443 11054
rect 15929 11051 15995 11054
rect 16205 11114 16271 11117
rect 16389 11114 16455 11117
rect 16205 11112 16455 11114
rect 16205 11056 16210 11112
rect 16266 11056 16394 11112
rect 16450 11056 16455 11112
rect 16205 11054 16455 11056
rect 16205 11051 16271 11054
rect 16389 11051 16455 11054
rect 15101 10980 15167 10981
rect 15101 10978 15148 10980
rect 15056 10976 15148 10978
rect 15056 10920 15106 10976
rect 15056 10918 15148 10920
rect 15101 10916 15148 10918
rect 15212 10916 15218 10980
rect 15101 10915 15167 10916
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 12606 10847 12922 10848
rect 17606 10912 17922 10913
rect 17606 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17922 10912
rect 17606 10847 17922 10848
rect 3785 10842 3851 10845
rect 3918 10842 3924 10844
rect 3785 10840 3924 10842
rect 3785 10784 3790 10840
rect 3846 10784 3924 10840
rect 3785 10782 3924 10784
rect 3785 10779 3851 10782
rect 3918 10780 3924 10782
rect 3988 10780 3994 10844
rect 11646 10780 11652 10844
rect 11716 10842 11722 10844
rect 11789 10842 11855 10845
rect 11716 10840 11855 10842
rect 11716 10784 11794 10840
rect 11850 10784 11855 10840
rect 11716 10782 11855 10784
rect 11716 10780 11722 10782
rect 11789 10779 11855 10782
rect 1209 10706 1275 10709
rect 13813 10706 13879 10709
rect 1209 10704 13879 10706
rect 1209 10648 1214 10704
rect 1270 10648 13818 10704
rect 13874 10648 13879 10704
rect 1209 10646 13879 10648
rect 1209 10643 1275 10646
rect 13813 10643 13879 10646
rect 6085 10570 6151 10573
rect 16481 10570 16547 10573
rect 6085 10568 16547 10570
rect 6085 10512 6090 10568
rect 6146 10512 16486 10568
rect 16542 10512 16547 10568
rect 6085 10510 16547 10512
rect 6085 10507 6151 10510
rect 16481 10507 16547 10510
rect 0 10434 800 10464
rect 0 10344 858 10434
rect 798 10301 858 10344
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 11946 10368 12262 10369
rect 11946 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12262 10368
rect 11946 10303 12262 10304
rect 16946 10368 17262 10369
rect 16946 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17262 10368
rect 16946 10303 17262 10304
rect 798 10296 907 10301
rect 798 10240 846 10296
rect 902 10240 907 10296
rect 798 10238 907 10240
rect 841 10235 907 10238
rect 7557 10298 7623 10301
rect 9070 10298 9076 10300
rect 7557 10296 9076 10298
rect 7557 10240 7562 10296
rect 7618 10240 9076 10296
rect 7557 10238 9076 10240
rect 7557 10235 7623 10238
rect 9070 10236 9076 10238
rect 9140 10298 9146 10300
rect 9622 10298 9628 10300
rect 9140 10238 9628 10298
rect 9140 10236 9146 10238
rect 9622 10236 9628 10238
rect 9692 10236 9698 10300
rect 12382 10236 12388 10300
rect 12452 10298 12458 10300
rect 15009 10298 15075 10301
rect 12452 10296 15075 10298
rect 12452 10240 15014 10296
rect 15070 10240 15075 10296
rect 12452 10238 15075 10240
rect 12452 10236 12458 10238
rect 15009 10235 15075 10238
rect 5073 10162 5139 10165
rect 9765 10162 9831 10165
rect 17861 10162 17927 10165
rect 5073 10160 9831 10162
rect 5073 10104 5078 10160
rect 5134 10104 9770 10160
rect 9826 10104 9831 10160
rect 5073 10102 9831 10104
rect 5073 10099 5139 10102
rect 9765 10099 9831 10102
rect 12344 10160 17927 10162
rect 12344 10104 17866 10160
rect 17922 10104 17927 10160
rect 12344 10102 17927 10104
rect 1393 10026 1459 10029
rect 2497 10026 2563 10029
rect 5533 10026 5599 10029
rect 12344 10026 12404 10102
rect 17861 10099 17927 10102
rect 1393 10024 5458 10026
rect 1393 9968 1398 10024
rect 1454 9968 2502 10024
rect 2558 9968 5458 10024
rect 1393 9966 5458 9968
rect 1393 9963 1459 9966
rect 2497 9963 2563 9966
rect 5398 9890 5458 9966
rect 5533 10024 12404 10026
rect 5533 9968 5538 10024
rect 5594 9968 12404 10024
rect 5533 9966 12404 9968
rect 16573 10026 16639 10029
rect 16798 10026 16804 10028
rect 16573 10024 16804 10026
rect 16573 9968 16578 10024
rect 16634 9968 16804 10024
rect 16573 9966 16804 9968
rect 5533 9963 5599 9966
rect 16573 9963 16639 9966
rect 16798 9964 16804 9966
rect 16868 9964 16874 10028
rect 8293 9890 8359 9893
rect 10542 9890 10548 9892
rect 5398 9830 7482 9890
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 3141 9754 3207 9757
rect 7281 9754 7347 9757
rect 3141 9752 7347 9754
rect 3141 9696 3146 9752
rect 3202 9696 7286 9752
rect 7342 9696 7347 9752
rect 3141 9694 7347 9696
rect 3141 9691 3207 9694
rect 7281 9691 7347 9694
rect 7422 9618 7482 9830
rect 8293 9888 10548 9890
rect 8293 9832 8298 9888
rect 8354 9832 10548 9888
rect 8293 9830 10548 9832
rect 8293 9827 8359 9830
rect 10542 9828 10548 9830
rect 10612 9890 10618 9892
rect 12382 9890 12388 9892
rect 10612 9830 12388 9890
rect 10612 9828 10618 9830
rect 12382 9828 12388 9830
rect 12452 9828 12458 9892
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 17606 9824 17922 9825
rect 17606 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17922 9824
rect 17606 9759 17922 9760
rect 10317 9754 10383 9757
rect 8158 9752 10383 9754
rect 8158 9696 10322 9752
rect 10378 9696 10383 9752
rect 8158 9694 10383 9696
rect 8158 9618 8218 9694
rect 10317 9691 10383 9694
rect 15193 9754 15259 9757
rect 15745 9754 15811 9757
rect 15193 9752 15811 9754
rect 15193 9696 15198 9752
rect 15254 9696 15750 9752
rect 15806 9696 15811 9752
rect 15193 9694 15811 9696
rect 15193 9691 15259 9694
rect 15745 9691 15811 9694
rect 7422 9558 8218 9618
rect 9581 9618 9647 9621
rect 16297 9618 16363 9621
rect 9581 9616 16363 9618
rect 9581 9560 9586 9616
rect 9642 9560 16302 9616
rect 16358 9560 16363 9616
rect 9581 9558 16363 9560
rect 9581 9555 9647 9558
rect 16297 9555 16363 9558
rect 841 9482 907 9485
rect 798 9480 907 9482
rect 798 9424 846 9480
rect 902 9424 907 9480
rect 798 9419 907 9424
rect 3693 9482 3759 9485
rect 6913 9482 6979 9485
rect 3693 9480 6979 9482
rect 3693 9424 3698 9480
rect 3754 9424 6918 9480
rect 6974 9424 6979 9480
rect 3693 9422 6979 9424
rect 3693 9419 3759 9422
rect 6913 9419 6979 9422
rect 11697 9482 11763 9485
rect 17125 9482 17191 9485
rect 11697 9480 17191 9482
rect 11697 9424 11702 9480
rect 11758 9424 17130 9480
rect 17186 9424 17191 9480
rect 11697 9422 17191 9424
rect 11697 9419 11763 9422
rect 17125 9419 17191 9422
rect 798 9376 858 9419
rect 0 9286 858 9376
rect 0 9256 800 9286
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 11946 9280 12262 9281
rect 11946 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12262 9280
rect 11946 9215 12262 9216
rect 16946 9280 17262 9281
rect 16946 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17262 9280
rect 16946 9215 17262 9216
rect 6545 9074 6611 9077
rect 17953 9074 18019 9077
rect 6545 9072 18019 9074
rect 6545 9016 6550 9072
rect 6606 9016 17958 9072
rect 18014 9016 18019 9072
rect 6545 9014 18019 9016
rect 6545 9011 6611 9014
rect 17953 9011 18019 9014
rect 2446 8876 2452 8940
rect 2516 8938 2522 8940
rect 2589 8938 2655 8941
rect 2516 8936 2655 8938
rect 2516 8880 2594 8936
rect 2650 8880 2655 8936
rect 2516 8878 2655 8880
rect 2516 8876 2522 8878
rect 2589 8875 2655 8878
rect 4061 8938 4127 8941
rect 13261 8938 13327 8941
rect 4061 8936 13327 8938
rect 4061 8880 4066 8936
rect 4122 8880 13266 8936
rect 13322 8880 13327 8936
rect 4061 8878 13327 8880
rect 4061 8875 4127 8878
rect 13261 8875 13327 8878
rect 14958 8876 14964 8940
rect 15028 8938 15034 8940
rect 15101 8938 15167 8941
rect 15028 8936 15167 8938
rect 15028 8880 15106 8936
rect 15162 8880 15167 8936
rect 15028 8878 15167 8880
rect 15028 8876 15034 8878
rect 15101 8875 15167 8878
rect 4061 8802 4127 8805
rect 6453 8802 6519 8805
rect 4061 8800 6519 8802
rect 4061 8744 4066 8800
rect 4122 8744 6458 8800
rect 6514 8744 6519 8800
rect 4061 8742 6519 8744
rect 4061 8739 4127 8742
rect 6453 8739 6519 8742
rect 8937 8802 9003 8805
rect 11697 8802 11763 8805
rect 8937 8800 11763 8802
rect 8937 8744 8942 8800
rect 8998 8744 11702 8800
rect 11758 8744 11763 8800
rect 8937 8742 11763 8744
rect 8937 8739 9003 8742
rect 11697 8739 11763 8742
rect 18413 8802 18479 8805
rect 19200 8802 20000 8832
rect 18413 8800 20000 8802
rect 18413 8744 18418 8800
rect 18474 8744 20000 8800
rect 18413 8742 20000 8744
rect 18413 8739 18479 8742
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 12606 8671 12922 8672
rect 17606 8736 17922 8737
rect 17606 8672 17612 8736
rect 17676 8672 17692 8736
rect 17756 8672 17772 8736
rect 17836 8672 17852 8736
rect 17916 8672 17922 8736
rect 19200 8712 20000 8742
rect 17606 8671 17922 8672
rect 13486 8530 13492 8532
rect 7790 8470 13492 8530
rect 3417 8394 3483 8397
rect 6637 8394 6703 8397
rect 3417 8392 6703 8394
rect 3417 8336 3422 8392
rect 3478 8336 6642 8392
rect 6698 8336 6703 8392
rect 3417 8334 6703 8336
rect 3417 8331 3483 8334
rect 6637 8331 6703 8334
rect 7414 8332 7420 8396
rect 7484 8394 7490 8396
rect 7649 8394 7715 8397
rect 7484 8392 7715 8394
rect 7484 8336 7654 8392
rect 7710 8336 7715 8392
rect 7484 8334 7715 8336
rect 7484 8332 7490 8334
rect 7649 8331 7715 8334
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 7373 8258 7439 8261
rect 7790 8258 7850 8470
rect 13486 8468 13492 8470
rect 13556 8530 13562 8532
rect 15193 8530 15259 8533
rect 13556 8528 15259 8530
rect 13556 8472 15198 8528
rect 15254 8472 15259 8528
rect 13556 8470 15259 8472
rect 13556 8468 13562 8470
rect 15193 8467 15259 8470
rect 9765 8394 9831 8397
rect 14089 8394 14155 8397
rect 9765 8392 14155 8394
rect 9765 8336 9770 8392
rect 9826 8336 14094 8392
rect 14150 8336 14155 8392
rect 9765 8334 14155 8336
rect 9765 8331 9831 8334
rect 14089 8331 14155 8334
rect 15377 8260 15443 8261
rect 15326 8258 15332 8260
rect 7373 8256 7850 8258
rect 7373 8200 7378 8256
rect 7434 8200 7850 8256
rect 7373 8198 7850 8200
rect 15286 8198 15332 8258
rect 15396 8256 15443 8260
rect 15438 8200 15443 8256
rect 7373 8195 7439 8198
rect 15326 8196 15332 8198
rect 15396 8196 15443 8200
rect 15377 8195 15443 8196
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 11946 8192 12262 8193
rect 11946 8128 11952 8192
rect 12016 8128 12032 8192
rect 12096 8128 12112 8192
rect 12176 8128 12192 8192
rect 12256 8128 12262 8192
rect 11946 8127 12262 8128
rect 16946 8192 17262 8193
rect 16946 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17262 8192
rect 16946 8127 17262 8128
rect 8109 8122 8175 8125
rect 8109 8120 8218 8122
rect 8109 8064 8114 8120
rect 8170 8064 8218 8120
rect 8109 8059 8218 8064
rect 8158 7986 8218 8059
rect 17677 7986 17743 7989
rect 8158 7984 17743 7986
rect 8158 7928 17682 7984
rect 17738 7928 17743 7984
rect 8158 7926 17743 7928
rect 17677 7923 17743 7926
rect 2313 7850 2379 7853
rect 3918 7850 3924 7852
rect 2313 7848 3924 7850
rect 2313 7792 2318 7848
rect 2374 7792 3924 7848
rect 2313 7790 3924 7792
rect 2313 7787 2379 7790
rect 3918 7788 3924 7790
rect 3988 7788 3994 7852
rect 7925 7850 7991 7853
rect 8150 7850 8156 7852
rect 7925 7848 8156 7850
rect 7925 7792 7930 7848
rect 7986 7792 8156 7848
rect 7925 7790 8156 7792
rect 7925 7787 7991 7790
rect 8150 7788 8156 7790
rect 8220 7788 8226 7852
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 12606 7583 12922 7584
rect 17606 7648 17922 7649
rect 17606 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17922 7648
rect 17606 7583 17922 7584
rect 841 7306 907 7309
rect 798 7304 907 7306
rect 798 7248 846 7304
rect 902 7248 907 7304
rect 798 7243 907 7248
rect 9806 7244 9812 7308
rect 9876 7306 9882 7308
rect 15653 7306 15719 7309
rect 9876 7304 15719 7306
rect 9876 7248 15658 7304
rect 15714 7248 15719 7304
rect 9876 7246 15719 7248
rect 9876 7244 9882 7246
rect 15653 7243 15719 7246
rect 798 7200 858 7243
rect 0 7110 858 7200
rect 0 7080 800 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 11946 7104 12262 7105
rect 11946 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12262 7104
rect 11946 7039 12262 7040
rect 16946 7104 17262 7105
rect 16946 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17262 7104
rect 16946 7039 17262 7040
rect 6126 6836 6132 6900
rect 6196 6898 6202 6900
rect 12525 6898 12591 6901
rect 6196 6896 12591 6898
rect 6196 6840 12530 6896
rect 12586 6840 12591 6896
rect 6196 6838 12591 6840
rect 6196 6836 6202 6838
rect 12525 6835 12591 6838
rect 13813 6898 13879 6901
rect 15101 6900 15167 6901
rect 14406 6898 14412 6900
rect 13813 6896 14412 6898
rect 13813 6840 13818 6896
rect 13874 6840 14412 6896
rect 13813 6838 14412 6840
rect 13813 6835 13879 6838
rect 14406 6836 14412 6838
rect 14476 6836 14482 6900
rect 15101 6896 15148 6900
rect 15212 6898 15218 6900
rect 15101 6840 15106 6896
rect 15101 6836 15148 6840
rect 15212 6838 15258 6898
rect 15212 6836 15218 6838
rect 15101 6835 15167 6836
rect 2037 6762 2103 6765
rect 4889 6762 4955 6765
rect 2037 6760 4955 6762
rect 2037 6704 2042 6760
rect 2098 6704 4894 6760
rect 4950 6704 4955 6760
rect 2037 6702 4955 6704
rect 2037 6699 2103 6702
rect 4889 6699 4955 6702
rect 8661 6762 8727 6765
rect 16113 6762 16179 6765
rect 8661 6760 16179 6762
rect 8661 6704 8666 6760
rect 8722 6704 16118 6760
rect 16174 6704 16179 6760
rect 8661 6702 16179 6704
rect 8661 6699 8727 6702
rect 16113 6699 16179 6702
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 12606 6495 12922 6496
rect 17606 6560 17922 6561
rect 17606 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17922 6560
rect 17606 6495 17922 6496
rect 13721 6492 13787 6493
rect 13670 6428 13676 6492
rect 13740 6490 13787 6492
rect 13740 6488 13832 6490
rect 13782 6432 13832 6488
rect 13740 6430 13832 6432
rect 13740 6428 13787 6430
rect 13721 6427 13787 6428
rect 8150 6292 8156 6356
rect 8220 6354 8226 6356
rect 18229 6354 18295 6357
rect 8220 6352 18295 6354
rect 8220 6296 18234 6352
rect 18290 6296 18295 6352
rect 8220 6294 18295 6296
rect 8220 6292 8226 6294
rect 18229 6291 18295 6294
rect 18413 6354 18479 6357
rect 19200 6354 20000 6384
rect 18413 6352 20000 6354
rect 18413 6296 18418 6352
rect 18474 6296 20000 6352
rect 18413 6294 20000 6296
rect 18413 6291 18479 6294
rect 19200 6264 20000 6294
rect 1761 6218 1827 6221
rect 14958 6218 14964 6220
rect 1761 6216 14964 6218
rect 1761 6160 1766 6216
rect 1822 6160 14964 6216
rect 1761 6158 14964 6160
rect 1761 6155 1827 6158
rect 14958 6156 14964 6158
rect 15028 6156 15034 6220
rect 0 6082 800 6112
rect 933 6082 999 6085
rect 0 6080 999 6082
rect 0 6024 938 6080
rect 994 6024 999 6080
rect 0 6022 999 6024
rect 0 5992 800 6022
rect 933 6019 999 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 11946 6016 12262 6017
rect 11946 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12262 6016
rect 11946 5951 12262 5952
rect 16946 6016 17262 6017
rect 16946 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17262 6016
rect 16946 5951 17262 5952
rect 13813 5946 13879 5949
rect 16757 5946 16823 5949
rect 7422 5886 11530 5946
rect 6729 5810 6795 5813
rect 7422 5810 7482 5886
rect 6729 5808 7482 5810
rect 6729 5752 6734 5808
rect 6790 5752 7482 5808
rect 6729 5750 7482 5752
rect 6729 5747 6795 5750
rect 9438 5748 9444 5812
rect 9508 5810 9514 5812
rect 11470 5810 11530 5886
rect 13813 5944 16823 5946
rect 13813 5888 13818 5944
rect 13874 5888 16762 5944
rect 16818 5888 16823 5944
rect 13813 5886 16823 5888
rect 13813 5883 13879 5886
rect 16757 5883 16823 5886
rect 14825 5810 14891 5813
rect 9508 5750 11300 5810
rect 11470 5808 14891 5810
rect 11470 5752 14830 5808
rect 14886 5752 14891 5808
rect 11470 5750 14891 5752
rect 9508 5748 9514 5750
rect 11094 5674 11100 5676
rect 9630 5614 11100 5674
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 3141 5266 3207 5269
rect 9630 5266 9690 5614
rect 11094 5612 11100 5614
rect 11164 5612 11170 5676
rect 11240 5538 11300 5750
rect 14825 5747 14891 5750
rect 11240 5478 12450 5538
rect 12249 5266 12315 5269
rect 3141 5264 9690 5266
rect 3141 5208 3146 5264
rect 3202 5208 9690 5264
rect 3141 5206 9690 5208
rect 10550 5264 12315 5266
rect 10550 5208 12254 5264
rect 12310 5208 12315 5264
rect 10550 5206 12315 5208
rect 12390 5266 12450 5478
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 12606 5407 12922 5408
rect 17606 5472 17922 5473
rect 17606 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17922 5472
rect 17606 5407 17922 5408
rect 14089 5266 14155 5269
rect 12390 5264 14155 5266
rect 12390 5208 14094 5264
rect 14150 5208 14155 5264
rect 12390 5206 14155 5208
rect 3141 5203 3207 5206
rect 841 5130 907 5133
rect 798 5128 907 5130
rect 798 5072 846 5128
rect 902 5072 907 5128
rect 798 5067 907 5072
rect 5165 5130 5231 5133
rect 8937 5130 9003 5133
rect 10550 5130 10610 5206
rect 12249 5203 12315 5206
rect 14089 5203 14155 5206
rect 5165 5128 7482 5130
rect 5165 5072 5170 5128
rect 5226 5072 7482 5128
rect 5165 5070 7482 5072
rect 5165 5067 5231 5070
rect 798 5024 858 5067
rect 0 4934 858 5024
rect 0 4904 800 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 7422 4858 7482 5070
rect 8937 5128 10610 5130
rect 8937 5072 8942 5128
rect 8998 5072 10610 5128
rect 8937 5070 10610 5072
rect 8937 5067 9003 5070
rect 10726 5068 10732 5132
rect 10796 5130 10802 5132
rect 13169 5130 13235 5133
rect 10796 5128 13235 5130
rect 10796 5072 13174 5128
rect 13230 5072 13235 5128
rect 10796 5070 13235 5072
rect 10796 5068 10802 5070
rect 13169 5067 13235 5070
rect 11946 4928 12262 4929
rect 11946 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12262 4928
rect 11946 4863 12262 4864
rect 16946 4928 17262 4929
rect 16946 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17262 4928
rect 16946 4863 17262 4864
rect 11145 4858 11211 4861
rect 11278 4858 11284 4860
rect 7422 4856 11284 4858
rect 7422 4800 11150 4856
rect 11206 4800 11284 4856
rect 7422 4798 11284 4800
rect 11145 4795 11211 4798
rect 11278 4796 11284 4798
rect 11348 4796 11354 4860
rect 6678 4660 6684 4724
rect 6748 4722 6754 4724
rect 12065 4722 12131 4725
rect 6748 4720 12131 4722
rect 6748 4664 12070 4720
rect 12126 4664 12131 4720
rect 6748 4662 12131 4664
rect 6748 4660 6754 4662
rect 12065 4659 12131 4662
rect 12249 4722 12315 4725
rect 15377 4722 15443 4725
rect 12249 4720 15443 4722
rect 12249 4664 12254 4720
rect 12310 4664 15382 4720
rect 15438 4664 15443 4720
rect 12249 4662 15443 4664
rect 12249 4659 12315 4662
rect 15377 4659 15443 4662
rect 2446 4524 2452 4588
rect 2516 4586 2522 4588
rect 15653 4586 15719 4589
rect 2516 4584 15719 4586
rect 2516 4528 15658 4584
rect 15714 4528 15719 4584
rect 2516 4526 15719 4528
rect 2516 4524 2522 4526
rect 15653 4523 15719 4526
rect 9029 4450 9095 4453
rect 12341 4450 12407 4453
rect 9029 4448 12407 4450
rect 9029 4392 9034 4448
rect 9090 4392 12346 4448
rect 12402 4392 12407 4448
rect 9029 4390 12407 4392
rect 9029 4387 9095 4390
rect 12341 4387 12407 4390
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 12606 4319 12922 4320
rect 17606 4384 17922 4385
rect 17606 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17922 4384
rect 17606 4319 17922 4320
rect 9806 4252 9812 4316
rect 9876 4314 9882 4316
rect 9949 4314 10015 4317
rect 9876 4312 10015 4314
rect 9876 4256 9954 4312
rect 10010 4256 10015 4312
rect 9876 4254 10015 4256
rect 9876 4252 9882 4254
rect 9949 4251 10015 4254
rect 6269 4178 6335 4181
rect 12249 4178 12315 4181
rect 6269 4176 12315 4178
rect 6269 4120 6274 4176
rect 6330 4120 12254 4176
rect 12310 4120 12315 4176
rect 6269 4118 12315 4120
rect 6269 4115 6335 4118
rect 12249 4115 12315 4118
rect 841 4042 907 4045
rect 798 4040 907 4042
rect 798 3984 846 4040
rect 902 3984 907 4040
rect 798 3979 907 3984
rect 5809 4042 5875 4045
rect 5942 4042 5948 4044
rect 5809 4040 5948 4042
rect 5809 3984 5814 4040
rect 5870 3984 5948 4040
rect 5809 3982 5948 3984
rect 5809 3979 5875 3982
rect 5942 3980 5948 3982
rect 6012 3980 6018 4044
rect 10133 4042 10199 4045
rect 12341 4042 12407 4045
rect 10133 4040 12407 4042
rect 10133 3984 10138 4040
rect 10194 3984 12346 4040
rect 12402 3984 12407 4040
rect 10133 3982 12407 3984
rect 10133 3979 10199 3982
rect 12341 3979 12407 3982
rect 798 3936 858 3979
rect 0 3846 858 3936
rect 18413 3906 18479 3909
rect 19200 3906 20000 3936
rect 18413 3904 20000 3906
rect 18413 3848 18418 3904
rect 18474 3848 20000 3904
rect 18413 3846 20000 3848
rect 0 3816 800 3846
rect 18413 3843 18479 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 11946 3840 12262 3841
rect 11946 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12262 3840
rect 11946 3775 12262 3776
rect 16946 3840 17262 3841
rect 16946 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17262 3840
rect 19200 3816 20000 3846
rect 16946 3775 17262 3776
rect 4654 3572 4660 3636
rect 4724 3634 4730 3636
rect 8845 3634 8911 3637
rect 4724 3632 8911 3634
rect 4724 3576 8850 3632
rect 8906 3576 8911 3632
rect 4724 3574 8911 3576
rect 4724 3572 4730 3574
rect 8845 3571 8911 3574
rect 5390 3436 5396 3500
rect 5460 3498 5466 3500
rect 14365 3498 14431 3501
rect 5460 3496 14431 3498
rect 5460 3440 14370 3496
rect 14426 3440 14431 3496
rect 5460 3438 14431 3440
rect 5460 3436 5466 3438
rect 14365 3435 14431 3438
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 12606 3231 12922 3232
rect 17606 3296 17922 3297
rect 17606 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17922 3296
rect 17606 3231 17922 3232
rect 10961 3228 11027 3229
rect 10910 3164 10916 3228
rect 10980 3226 11027 3228
rect 10980 3224 11072 3226
rect 11022 3168 11072 3224
rect 10980 3166 11072 3168
rect 10980 3164 11027 3166
rect 10961 3163 11027 3164
rect 841 2954 907 2957
rect 798 2952 907 2954
rect 798 2896 846 2952
rect 902 2896 907 2952
rect 798 2891 907 2896
rect 2313 2954 2379 2957
rect 16614 2954 16620 2956
rect 2313 2952 16620 2954
rect 2313 2896 2318 2952
rect 2374 2896 16620 2952
rect 2313 2894 16620 2896
rect 2313 2891 2379 2894
rect 16614 2892 16620 2894
rect 16684 2892 16690 2956
rect 798 2848 858 2891
rect 0 2758 858 2848
rect 0 2728 800 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 11946 2752 12262 2753
rect 11946 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12262 2752
rect 11946 2687 12262 2688
rect 16946 2752 17262 2753
rect 16946 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17262 2752
rect 16946 2687 17262 2688
rect 9121 2682 9187 2685
rect 9254 2682 9260 2684
rect 9121 2680 9260 2682
rect 9121 2624 9126 2680
rect 9182 2624 9260 2680
rect 9121 2622 9260 2624
rect 9121 2619 9187 2622
rect 9254 2620 9260 2622
rect 9324 2620 9330 2684
rect 15745 2546 15811 2549
rect 15878 2546 15884 2548
rect 15745 2544 15884 2546
rect 15745 2488 15750 2544
rect 15806 2488 15884 2544
rect 15745 2486 15884 2488
rect 15745 2483 15811 2486
rect 15878 2484 15884 2486
rect 15948 2484 15954 2548
rect 6494 2348 6500 2412
rect 6564 2410 6570 2412
rect 16113 2410 16179 2413
rect 6564 2408 16179 2410
rect 6564 2352 16118 2408
rect 16174 2352 16179 2408
rect 6564 2350 16179 2352
rect 6564 2348 6570 2350
rect 16113 2347 16179 2350
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 12606 2143 12922 2144
rect 17606 2208 17922 2209
rect 17606 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17922 2208
rect 17606 2143 17922 2144
rect 0 1730 800 1760
rect 1853 1730 1919 1733
rect 0 1728 1919 1730
rect 0 1672 1858 1728
rect 1914 1672 1919 1728
rect 0 1670 1919 1672
rect 0 1640 800 1670
rect 1853 1667 1919 1670
rect 18413 1458 18479 1461
rect 19200 1458 20000 1488
rect 18413 1456 20000 1458
rect 18413 1400 18418 1456
rect 18474 1400 20000 1456
rect 18413 1398 20000 1400
rect 18413 1395 18479 1398
rect 19200 1368 20000 1398
<< via3 >>
rect 2612 17436 2676 17440
rect 2612 17380 2616 17436
rect 2616 17380 2672 17436
rect 2672 17380 2676 17436
rect 2612 17376 2676 17380
rect 2692 17436 2756 17440
rect 2692 17380 2696 17436
rect 2696 17380 2752 17436
rect 2752 17380 2756 17436
rect 2692 17376 2756 17380
rect 2772 17436 2836 17440
rect 2772 17380 2776 17436
rect 2776 17380 2832 17436
rect 2832 17380 2836 17436
rect 2772 17376 2836 17380
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 7612 17436 7676 17440
rect 7612 17380 7616 17436
rect 7616 17380 7672 17436
rect 7672 17380 7676 17436
rect 7612 17376 7676 17380
rect 7692 17436 7756 17440
rect 7692 17380 7696 17436
rect 7696 17380 7752 17436
rect 7752 17380 7756 17436
rect 7692 17376 7756 17380
rect 7772 17436 7836 17440
rect 7772 17380 7776 17436
rect 7776 17380 7832 17436
rect 7832 17380 7836 17436
rect 7772 17376 7836 17380
rect 7852 17436 7916 17440
rect 7852 17380 7856 17436
rect 7856 17380 7912 17436
rect 7912 17380 7916 17436
rect 7852 17376 7916 17380
rect 12612 17436 12676 17440
rect 12612 17380 12616 17436
rect 12616 17380 12672 17436
rect 12672 17380 12676 17436
rect 12612 17376 12676 17380
rect 12692 17436 12756 17440
rect 12692 17380 12696 17436
rect 12696 17380 12752 17436
rect 12752 17380 12756 17436
rect 12692 17376 12756 17380
rect 12772 17436 12836 17440
rect 12772 17380 12776 17436
rect 12776 17380 12832 17436
rect 12832 17380 12836 17436
rect 12772 17376 12836 17380
rect 12852 17436 12916 17440
rect 12852 17380 12856 17436
rect 12856 17380 12912 17436
rect 12912 17380 12916 17436
rect 12852 17376 12916 17380
rect 17612 17436 17676 17440
rect 17612 17380 17616 17436
rect 17616 17380 17672 17436
rect 17672 17380 17676 17436
rect 17612 17376 17676 17380
rect 17692 17436 17756 17440
rect 17692 17380 17696 17436
rect 17696 17380 17752 17436
rect 17752 17380 17756 17436
rect 17692 17376 17756 17380
rect 17772 17436 17836 17440
rect 17772 17380 17776 17436
rect 17776 17380 17832 17436
rect 17832 17380 17836 17436
rect 17772 17376 17836 17380
rect 17852 17436 17916 17440
rect 17852 17380 17856 17436
rect 17856 17380 17912 17436
rect 17912 17380 17916 17436
rect 17852 17376 17916 17380
rect 5948 17036 6012 17100
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 6952 16892 7016 16896
rect 6952 16836 6956 16892
rect 6956 16836 7012 16892
rect 7012 16836 7016 16892
rect 6952 16832 7016 16836
rect 7032 16892 7096 16896
rect 7032 16836 7036 16892
rect 7036 16836 7092 16892
rect 7092 16836 7096 16892
rect 7032 16832 7096 16836
rect 7112 16892 7176 16896
rect 7112 16836 7116 16892
rect 7116 16836 7172 16892
rect 7172 16836 7176 16892
rect 7112 16832 7176 16836
rect 7192 16892 7256 16896
rect 7192 16836 7196 16892
rect 7196 16836 7252 16892
rect 7252 16836 7256 16892
rect 7192 16832 7256 16836
rect 11952 16892 12016 16896
rect 11952 16836 11956 16892
rect 11956 16836 12012 16892
rect 12012 16836 12016 16892
rect 11952 16832 12016 16836
rect 12032 16892 12096 16896
rect 12032 16836 12036 16892
rect 12036 16836 12092 16892
rect 12092 16836 12096 16892
rect 12032 16832 12096 16836
rect 12112 16892 12176 16896
rect 12112 16836 12116 16892
rect 12116 16836 12172 16892
rect 12172 16836 12176 16892
rect 12112 16832 12176 16836
rect 12192 16892 12256 16896
rect 12192 16836 12196 16892
rect 12196 16836 12252 16892
rect 12252 16836 12256 16892
rect 12192 16832 12256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 11100 16628 11164 16692
rect 14412 16356 14476 16420
rect 2612 16348 2676 16352
rect 2612 16292 2616 16348
rect 2616 16292 2672 16348
rect 2672 16292 2676 16348
rect 2612 16288 2676 16292
rect 2692 16348 2756 16352
rect 2692 16292 2696 16348
rect 2696 16292 2752 16348
rect 2752 16292 2756 16348
rect 2692 16288 2756 16292
rect 2772 16348 2836 16352
rect 2772 16292 2776 16348
rect 2776 16292 2832 16348
rect 2832 16292 2836 16348
rect 2772 16288 2836 16292
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 7612 16348 7676 16352
rect 7612 16292 7616 16348
rect 7616 16292 7672 16348
rect 7672 16292 7676 16348
rect 7612 16288 7676 16292
rect 7692 16348 7756 16352
rect 7692 16292 7696 16348
rect 7696 16292 7752 16348
rect 7752 16292 7756 16348
rect 7692 16288 7756 16292
rect 7772 16348 7836 16352
rect 7772 16292 7776 16348
rect 7776 16292 7832 16348
rect 7832 16292 7836 16348
rect 7772 16288 7836 16292
rect 7852 16348 7916 16352
rect 7852 16292 7856 16348
rect 7856 16292 7912 16348
rect 7912 16292 7916 16348
rect 7852 16288 7916 16292
rect 12612 16348 12676 16352
rect 12612 16292 12616 16348
rect 12616 16292 12672 16348
rect 12672 16292 12676 16348
rect 12612 16288 12676 16292
rect 12692 16348 12756 16352
rect 12692 16292 12696 16348
rect 12696 16292 12752 16348
rect 12752 16292 12756 16348
rect 12692 16288 12756 16292
rect 12772 16348 12836 16352
rect 12772 16292 12776 16348
rect 12776 16292 12832 16348
rect 12832 16292 12836 16348
rect 12772 16288 12836 16292
rect 12852 16348 12916 16352
rect 12852 16292 12856 16348
rect 12856 16292 12912 16348
rect 12912 16292 12916 16348
rect 12852 16288 12916 16292
rect 17612 16348 17676 16352
rect 17612 16292 17616 16348
rect 17616 16292 17672 16348
rect 17672 16292 17676 16348
rect 17612 16288 17676 16292
rect 17692 16348 17756 16352
rect 17692 16292 17696 16348
rect 17696 16292 17752 16348
rect 17752 16292 17756 16348
rect 17692 16288 17756 16292
rect 17772 16348 17836 16352
rect 17772 16292 17776 16348
rect 17776 16292 17832 16348
rect 17832 16292 17836 16348
rect 17772 16288 17836 16292
rect 17852 16348 17916 16352
rect 17852 16292 17856 16348
rect 17856 16292 17912 16348
rect 17912 16292 17916 16348
rect 17852 16288 17916 16292
rect 4660 15948 4724 16012
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 6952 15804 7016 15808
rect 6952 15748 6956 15804
rect 6956 15748 7012 15804
rect 7012 15748 7016 15804
rect 6952 15744 7016 15748
rect 7032 15804 7096 15808
rect 7032 15748 7036 15804
rect 7036 15748 7092 15804
rect 7092 15748 7096 15804
rect 7032 15744 7096 15748
rect 7112 15804 7176 15808
rect 7112 15748 7116 15804
rect 7116 15748 7172 15804
rect 7172 15748 7176 15804
rect 7112 15744 7176 15748
rect 7192 15804 7256 15808
rect 7192 15748 7196 15804
rect 7196 15748 7252 15804
rect 7252 15748 7256 15804
rect 7192 15744 7256 15748
rect 11952 15804 12016 15808
rect 11952 15748 11956 15804
rect 11956 15748 12012 15804
rect 12012 15748 12016 15804
rect 11952 15744 12016 15748
rect 12032 15804 12096 15808
rect 12032 15748 12036 15804
rect 12036 15748 12092 15804
rect 12092 15748 12096 15804
rect 12032 15744 12096 15748
rect 12112 15804 12176 15808
rect 12112 15748 12116 15804
rect 12116 15748 12172 15804
rect 12172 15748 12176 15804
rect 12112 15744 12176 15748
rect 12192 15804 12256 15808
rect 12192 15748 12196 15804
rect 12196 15748 12252 15804
rect 12252 15748 12256 15804
rect 12192 15744 12256 15748
rect 9260 15540 9324 15604
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 16620 15540 16684 15604
rect 6500 15404 6564 15468
rect 6684 15328 6748 15332
rect 6684 15272 6698 15328
rect 6698 15272 6748 15328
rect 6684 15268 6748 15272
rect 9444 15328 9508 15332
rect 9444 15272 9458 15328
rect 9458 15272 9508 15328
rect 9444 15268 9508 15272
rect 10364 15328 10428 15332
rect 10364 15272 10414 15328
rect 10414 15272 10428 15328
rect 10364 15268 10428 15272
rect 10732 15268 10796 15332
rect 10916 15328 10980 15332
rect 10916 15272 10966 15328
rect 10966 15272 10980 15328
rect 10916 15268 10980 15272
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 7612 15260 7676 15264
rect 7612 15204 7616 15260
rect 7616 15204 7672 15260
rect 7672 15204 7676 15260
rect 7612 15200 7676 15204
rect 7692 15260 7756 15264
rect 7692 15204 7696 15260
rect 7696 15204 7752 15260
rect 7752 15204 7756 15260
rect 7692 15200 7756 15204
rect 7772 15260 7836 15264
rect 7772 15204 7776 15260
rect 7776 15204 7832 15260
rect 7832 15204 7836 15260
rect 7772 15200 7836 15204
rect 7852 15260 7916 15264
rect 7852 15204 7856 15260
rect 7856 15204 7912 15260
rect 7912 15204 7916 15260
rect 7852 15200 7916 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 17612 15260 17676 15264
rect 17612 15204 17616 15260
rect 17616 15204 17672 15260
rect 17672 15204 17676 15260
rect 17612 15200 17676 15204
rect 17692 15260 17756 15264
rect 17692 15204 17696 15260
rect 17696 15204 17752 15260
rect 17752 15204 17756 15260
rect 17692 15200 17756 15204
rect 17772 15260 17836 15264
rect 17772 15204 17776 15260
rect 17776 15204 17832 15260
rect 17832 15204 17836 15260
rect 17772 15200 17836 15204
rect 17852 15260 17916 15264
rect 17852 15204 17856 15260
rect 17856 15204 17912 15260
rect 17912 15204 17916 15260
rect 17852 15200 17916 15204
rect 9812 14724 9876 14788
rect 10548 14784 10612 14788
rect 10548 14728 10598 14784
rect 10598 14728 10612 14784
rect 10548 14724 10612 14728
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 6952 14716 7016 14720
rect 6952 14660 6956 14716
rect 6956 14660 7012 14716
rect 7012 14660 7016 14716
rect 6952 14656 7016 14660
rect 7032 14716 7096 14720
rect 7032 14660 7036 14716
rect 7036 14660 7092 14716
rect 7092 14660 7096 14716
rect 7032 14656 7096 14660
rect 7112 14716 7176 14720
rect 7112 14660 7116 14716
rect 7116 14660 7172 14716
rect 7172 14660 7176 14716
rect 7112 14656 7176 14660
rect 7192 14716 7256 14720
rect 7192 14660 7196 14716
rect 7196 14660 7252 14716
rect 7252 14660 7256 14716
rect 7192 14656 7256 14660
rect 11952 14716 12016 14720
rect 11952 14660 11956 14716
rect 11956 14660 12012 14716
rect 12012 14660 12016 14716
rect 11952 14656 12016 14660
rect 12032 14716 12096 14720
rect 12032 14660 12036 14716
rect 12036 14660 12092 14716
rect 12092 14660 12096 14716
rect 12032 14656 12096 14660
rect 12112 14716 12176 14720
rect 12112 14660 12116 14716
rect 12116 14660 12172 14716
rect 12172 14660 12176 14716
rect 12112 14656 12176 14660
rect 12192 14716 12256 14720
rect 12192 14660 12196 14716
rect 12196 14660 12252 14716
rect 12252 14660 12256 14716
rect 12192 14656 12256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 9996 14452 10060 14516
rect 3924 14316 3988 14380
rect 15332 14316 15396 14380
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 7612 14172 7676 14176
rect 7612 14116 7616 14172
rect 7616 14116 7672 14172
rect 7672 14116 7676 14172
rect 7612 14112 7676 14116
rect 7692 14172 7756 14176
rect 7692 14116 7696 14172
rect 7696 14116 7752 14172
rect 7752 14116 7756 14172
rect 7692 14112 7756 14116
rect 7772 14172 7836 14176
rect 7772 14116 7776 14172
rect 7776 14116 7832 14172
rect 7832 14116 7836 14172
rect 7772 14112 7836 14116
rect 7852 14172 7916 14176
rect 7852 14116 7856 14172
rect 7856 14116 7912 14172
rect 7912 14116 7916 14172
rect 7852 14112 7916 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 17612 14172 17676 14176
rect 17612 14116 17616 14172
rect 17616 14116 17672 14172
rect 17672 14116 17676 14172
rect 17612 14112 17676 14116
rect 17692 14172 17756 14176
rect 17692 14116 17696 14172
rect 17696 14116 17752 14172
rect 17752 14116 17756 14172
rect 17692 14112 17756 14116
rect 17772 14172 17836 14176
rect 17772 14116 17776 14172
rect 17776 14116 17832 14172
rect 17832 14116 17836 14172
rect 17772 14112 17836 14116
rect 17852 14172 17916 14176
rect 17852 14116 17856 14172
rect 17856 14116 17912 14172
rect 17912 14116 17916 14172
rect 17852 14112 17916 14116
rect 8156 13908 8220 13972
rect 6132 13772 6196 13836
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 6952 13628 7016 13632
rect 6952 13572 6956 13628
rect 6956 13572 7012 13628
rect 7012 13572 7016 13628
rect 6952 13568 7016 13572
rect 7032 13628 7096 13632
rect 7032 13572 7036 13628
rect 7036 13572 7092 13628
rect 7092 13572 7096 13628
rect 7032 13568 7096 13572
rect 7112 13628 7176 13632
rect 7112 13572 7116 13628
rect 7116 13572 7172 13628
rect 7172 13572 7176 13628
rect 7112 13568 7176 13572
rect 7192 13628 7256 13632
rect 7192 13572 7196 13628
rect 7196 13572 7252 13628
rect 7252 13572 7256 13628
rect 7192 13568 7256 13572
rect 9076 13500 9140 13564
rect 13492 13772 13556 13836
rect 14964 13772 15028 13836
rect 11952 13628 12016 13632
rect 11952 13572 11956 13628
rect 11956 13572 12012 13628
rect 12012 13572 12016 13628
rect 11952 13568 12016 13572
rect 12032 13628 12096 13632
rect 12032 13572 12036 13628
rect 12036 13572 12092 13628
rect 12092 13572 12096 13628
rect 12032 13568 12096 13572
rect 12112 13628 12176 13632
rect 12112 13572 12116 13628
rect 12116 13572 12172 13628
rect 12172 13572 12176 13628
rect 12112 13568 12176 13572
rect 12192 13628 12256 13632
rect 12192 13572 12196 13628
rect 12196 13572 12252 13628
rect 12252 13572 12256 13628
rect 12192 13568 12256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 15884 13500 15948 13564
rect 7420 13228 7484 13292
rect 13676 13364 13740 13428
rect 9260 13092 9324 13156
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 7612 13084 7676 13088
rect 7612 13028 7616 13084
rect 7616 13028 7672 13084
rect 7672 13028 7676 13084
rect 7612 13024 7676 13028
rect 7692 13084 7756 13088
rect 7692 13028 7696 13084
rect 7696 13028 7752 13084
rect 7752 13028 7756 13084
rect 7692 13024 7756 13028
rect 7772 13084 7836 13088
rect 7772 13028 7776 13084
rect 7776 13028 7832 13084
rect 7832 13028 7836 13084
rect 7772 13024 7836 13028
rect 7852 13084 7916 13088
rect 7852 13028 7856 13084
rect 7856 13028 7912 13084
rect 7912 13028 7916 13084
rect 7852 13024 7916 13028
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 17612 13084 17676 13088
rect 17612 13028 17616 13084
rect 17616 13028 17672 13084
rect 17672 13028 17676 13084
rect 17612 13024 17676 13028
rect 17692 13084 17756 13088
rect 17692 13028 17696 13084
rect 17696 13028 17752 13084
rect 17752 13028 17756 13084
rect 17692 13024 17756 13028
rect 17772 13084 17836 13088
rect 17772 13028 17776 13084
rect 17776 13028 17832 13084
rect 17832 13028 17836 13084
rect 17772 13024 17836 13028
rect 17852 13084 17916 13088
rect 17852 13028 17856 13084
rect 17856 13028 17912 13084
rect 17912 13028 17916 13084
rect 17852 13024 17916 13028
rect 5396 12684 5460 12748
rect 16804 12744 16868 12748
rect 16804 12688 16854 12744
rect 16854 12688 16868 12744
rect 16804 12684 16868 12688
rect 17356 12744 17420 12748
rect 17356 12688 17370 12744
rect 17370 12688 17420 12744
rect 17356 12684 17420 12688
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 6952 12540 7016 12544
rect 6952 12484 6956 12540
rect 6956 12484 7012 12540
rect 7012 12484 7016 12540
rect 6952 12480 7016 12484
rect 7032 12540 7096 12544
rect 7032 12484 7036 12540
rect 7036 12484 7092 12540
rect 7092 12484 7096 12540
rect 7032 12480 7096 12484
rect 7112 12540 7176 12544
rect 7112 12484 7116 12540
rect 7116 12484 7172 12540
rect 7172 12484 7176 12540
rect 7112 12480 7176 12484
rect 7192 12540 7256 12544
rect 7192 12484 7196 12540
rect 7196 12484 7252 12540
rect 7252 12484 7256 12540
rect 7192 12480 7256 12484
rect 11952 12540 12016 12544
rect 11952 12484 11956 12540
rect 11956 12484 12012 12540
rect 12012 12484 12016 12540
rect 11952 12480 12016 12484
rect 12032 12540 12096 12544
rect 12032 12484 12036 12540
rect 12036 12484 12092 12540
rect 12092 12484 12096 12540
rect 12032 12480 12096 12484
rect 12112 12540 12176 12544
rect 12112 12484 12116 12540
rect 12116 12484 12172 12540
rect 12172 12484 12176 12540
rect 12112 12480 12176 12484
rect 12192 12540 12256 12544
rect 12192 12484 12196 12540
rect 12196 12484 12252 12540
rect 12252 12484 12256 12540
rect 12192 12480 12256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 8156 12276 8220 12340
rect 17356 12336 17420 12340
rect 17356 12280 17406 12336
rect 17406 12280 17420 12336
rect 17356 12276 17420 12280
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 7612 11996 7676 12000
rect 7612 11940 7616 11996
rect 7616 11940 7672 11996
rect 7672 11940 7676 11996
rect 7612 11936 7676 11940
rect 7692 11996 7756 12000
rect 7692 11940 7696 11996
rect 7696 11940 7752 11996
rect 7752 11940 7756 11996
rect 7692 11936 7756 11940
rect 7772 11996 7836 12000
rect 7772 11940 7776 11996
rect 7776 11940 7832 11996
rect 7832 11940 7836 11996
rect 7772 11936 7836 11940
rect 7852 11996 7916 12000
rect 7852 11940 7856 11996
rect 7856 11940 7912 11996
rect 7912 11940 7916 11996
rect 7852 11936 7916 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 17612 11996 17676 12000
rect 17612 11940 17616 11996
rect 17616 11940 17672 11996
rect 17672 11940 17676 11996
rect 17612 11936 17676 11940
rect 17692 11996 17756 12000
rect 17692 11940 17696 11996
rect 17696 11940 17752 11996
rect 17752 11940 17756 11996
rect 17692 11936 17756 11940
rect 17772 11996 17836 12000
rect 17772 11940 17776 11996
rect 17776 11940 17832 11996
rect 17832 11940 17836 11996
rect 17772 11936 17836 11940
rect 17852 11996 17916 12000
rect 17852 11940 17856 11996
rect 17856 11940 17912 11996
rect 17912 11940 17916 11996
rect 17852 11936 17916 11940
rect 10364 11868 10428 11932
rect 11652 11868 11716 11932
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 11952 11452 12016 11456
rect 11952 11396 11956 11452
rect 11956 11396 12012 11452
rect 12012 11396 12016 11452
rect 11952 11392 12016 11396
rect 12032 11452 12096 11456
rect 12032 11396 12036 11452
rect 12036 11396 12092 11452
rect 12092 11396 12096 11452
rect 12032 11392 12096 11396
rect 12112 11452 12176 11456
rect 12112 11396 12116 11452
rect 12116 11396 12172 11452
rect 12172 11396 12176 11452
rect 12112 11392 12176 11396
rect 12192 11452 12256 11456
rect 12192 11396 12196 11452
rect 12196 11396 12252 11452
rect 12252 11396 12256 11452
rect 12192 11392 12256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 11100 11324 11164 11388
rect 15148 10976 15212 10980
rect 15148 10920 15162 10976
rect 15162 10920 15212 10976
rect 15148 10916 15212 10920
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 17612 10908 17676 10912
rect 17612 10852 17616 10908
rect 17616 10852 17672 10908
rect 17672 10852 17676 10908
rect 17612 10848 17676 10852
rect 17692 10908 17756 10912
rect 17692 10852 17696 10908
rect 17696 10852 17752 10908
rect 17752 10852 17756 10908
rect 17692 10848 17756 10852
rect 17772 10908 17836 10912
rect 17772 10852 17776 10908
rect 17776 10852 17832 10908
rect 17832 10852 17836 10908
rect 17772 10848 17836 10852
rect 17852 10908 17916 10912
rect 17852 10852 17856 10908
rect 17856 10852 17912 10908
rect 17912 10852 17916 10908
rect 17852 10848 17916 10852
rect 3924 10780 3988 10844
rect 11652 10780 11716 10844
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 11952 10364 12016 10368
rect 11952 10308 11956 10364
rect 11956 10308 12012 10364
rect 12012 10308 12016 10364
rect 11952 10304 12016 10308
rect 12032 10364 12096 10368
rect 12032 10308 12036 10364
rect 12036 10308 12092 10364
rect 12092 10308 12096 10364
rect 12032 10304 12096 10308
rect 12112 10364 12176 10368
rect 12112 10308 12116 10364
rect 12116 10308 12172 10364
rect 12172 10308 12176 10364
rect 12112 10304 12176 10308
rect 12192 10364 12256 10368
rect 12192 10308 12196 10364
rect 12196 10308 12252 10364
rect 12252 10308 12256 10364
rect 12192 10304 12256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 9076 10236 9140 10300
rect 9628 10236 9692 10300
rect 12388 10236 12452 10300
rect 16804 9964 16868 10028
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 10548 9828 10612 9892
rect 12388 9828 12452 9892
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 17612 9820 17676 9824
rect 17612 9764 17616 9820
rect 17616 9764 17672 9820
rect 17672 9764 17676 9820
rect 17612 9760 17676 9764
rect 17692 9820 17756 9824
rect 17692 9764 17696 9820
rect 17696 9764 17752 9820
rect 17752 9764 17756 9820
rect 17692 9760 17756 9764
rect 17772 9820 17836 9824
rect 17772 9764 17776 9820
rect 17776 9764 17832 9820
rect 17832 9764 17836 9820
rect 17772 9760 17836 9764
rect 17852 9820 17916 9824
rect 17852 9764 17856 9820
rect 17856 9764 17912 9820
rect 17912 9764 17916 9820
rect 17852 9760 17916 9764
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 11952 9276 12016 9280
rect 11952 9220 11956 9276
rect 11956 9220 12012 9276
rect 12012 9220 12016 9276
rect 11952 9216 12016 9220
rect 12032 9276 12096 9280
rect 12032 9220 12036 9276
rect 12036 9220 12092 9276
rect 12092 9220 12096 9276
rect 12032 9216 12096 9220
rect 12112 9276 12176 9280
rect 12112 9220 12116 9276
rect 12116 9220 12172 9276
rect 12172 9220 12176 9276
rect 12112 9216 12176 9220
rect 12192 9276 12256 9280
rect 12192 9220 12196 9276
rect 12196 9220 12252 9276
rect 12252 9220 12256 9276
rect 12192 9216 12256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 2452 8876 2516 8940
rect 14964 8876 15028 8940
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 17612 8732 17676 8736
rect 17612 8676 17616 8732
rect 17616 8676 17672 8732
rect 17672 8676 17676 8732
rect 17612 8672 17676 8676
rect 17692 8732 17756 8736
rect 17692 8676 17696 8732
rect 17696 8676 17752 8732
rect 17752 8676 17756 8732
rect 17692 8672 17756 8676
rect 17772 8732 17836 8736
rect 17772 8676 17776 8732
rect 17776 8676 17832 8732
rect 17832 8676 17836 8732
rect 17772 8672 17836 8676
rect 17852 8732 17916 8736
rect 17852 8676 17856 8732
rect 17856 8676 17912 8732
rect 17912 8676 17916 8732
rect 17852 8672 17916 8676
rect 7420 8332 7484 8396
rect 13492 8468 13556 8532
rect 15332 8256 15396 8260
rect 15332 8200 15382 8256
rect 15382 8200 15396 8256
rect 15332 8196 15396 8200
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 11952 8188 12016 8192
rect 11952 8132 11956 8188
rect 11956 8132 12012 8188
rect 12012 8132 12016 8188
rect 11952 8128 12016 8132
rect 12032 8188 12096 8192
rect 12032 8132 12036 8188
rect 12036 8132 12092 8188
rect 12092 8132 12096 8188
rect 12032 8128 12096 8132
rect 12112 8188 12176 8192
rect 12112 8132 12116 8188
rect 12116 8132 12172 8188
rect 12172 8132 12176 8188
rect 12112 8128 12176 8132
rect 12192 8188 12256 8192
rect 12192 8132 12196 8188
rect 12196 8132 12252 8188
rect 12252 8132 12256 8188
rect 12192 8128 12256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 3924 7788 3988 7852
rect 8156 7788 8220 7852
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 17612 7644 17676 7648
rect 17612 7588 17616 7644
rect 17616 7588 17672 7644
rect 17672 7588 17676 7644
rect 17612 7584 17676 7588
rect 17692 7644 17756 7648
rect 17692 7588 17696 7644
rect 17696 7588 17752 7644
rect 17752 7588 17756 7644
rect 17692 7584 17756 7588
rect 17772 7644 17836 7648
rect 17772 7588 17776 7644
rect 17776 7588 17832 7644
rect 17832 7588 17836 7644
rect 17772 7584 17836 7588
rect 17852 7644 17916 7648
rect 17852 7588 17856 7644
rect 17856 7588 17912 7644
rect 17912 7588 17916 7644
rect 17852 7584 17916 7588
rect 9812 7244 9876 7308
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 11952 7100 12016 7104
rect 11952 7044 11956 7100
rect 11956 7044 12012 7100
rect 12012 7044 12016 7100
rect 11952 7040 12016 7044
rect 12032 7100 12096 7104
rect 12032 7044 12036 7100
rect 12036 7044 12092 7100
rect 12092 7044 12096 7100
rect 12032 7040 12096 7044
rect 12112 7100 12176 7104
rect 12112 7044 12116 7100
rect 12116 7044 12172 7100
rect 12172 7044 12176 7100
rect 12112 7040 12176 7044
rect 12192 7100 12256 7104
rect 12192 7044 12196 7100
rect 12196 7044 12252 7100
rect 12252 7044 12256 7100
rect 12192 7040 12256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 6132 6836 6196 6900
rect 14412 6836 14476 6900
rect 15148 6896 15212 6900
rect 15148 6840 15162 6896
rect 15162 6840 15212 6896
rect 15148 6836 15212 6840
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 17612 6556 17676 6560
rect 17612 6500 17616 6556
rect 17616 6500 17672 6556
rect 17672 6500 17676 6556
rect 17612 6496 17676 6500
rect 17692 6556 17756 6560
rect 17692 6500 17696 6556
rect 17696 6500 17752 6556
rect 17752 6500 17756 6556
rect 17692 6496 17756 6500
rect 17772 6556 17836 6560
rect 17772 6500 17776 6556
rect 17776 6500 17832 6556
rect 17832 6500 17836 6556
rect 17772 6496 17836 6500
rect 17852 6556 17916 6560
rect 17852 6500 17856 6556
rect 17856 6500 17912 6556
rect 17912 6500 17916 6556
rect 17852 6496 17916 6500
rect 13676 6488 13740 6492
rect 13676 6432 13726 6488
rect 13726 6432 13740 6488
rect 13676 6428 13740 6432
rect 8156 6292 8220 6356
rect 14964 6156 15028 6220
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 11952 6012 12016 6016
rect 11952 5956 11956 6012
rect 11956 5956 12012 6012
rect 12012 5956 12016 6012
rect 11952 5952 12016 5956
rect 12032 6012 12096 6016
rect 12032 5956 12036 6012
rect 12036 5956 12092 6012
rect 12092 5956 12096 6012
rect 12032 5952 12096 5956
rect 12112 6012 12176 6016
rect 12112 5956 12116 6012
rect 12116 5956 12172 6012
rect 12172 5956 12176 6012
rect 12112 5952 12176 5956
rect 12192 6012 12256 6016
rect 12192 5956 12196 6012
rect 12196 5956 12252 6012
rect 12252 5956 12256 6012
rect 12192 5952 12256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 9444 5748 9508 5812
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 11100 5612 11164 5676
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 17612 5468 17676 5472
rect 17612 5412 17616 5468
rect 17616 5412 17672 5468
rect 17672 5412 17676 5468
rect 17612 5408 17676 5412
rect 17692 5468 17756 5472
rect 17692 5412 17696 5468
rect 17696 5412 17752 5468
rect 17752 5412 17756 5468
rect 17692 5408 17756 5412
rect 17772 5468 17836 5472
rect 17772 5412 17776 5468
rect 17776 5412 17832 5468
rect 17832 5412 17836 5468
rect 17772 5408 17836 5412
rect 17852 5468 17916 5472
rect 17852 5412 17856 5468
rect 17856 5412 17912 5468
rect 17912 5412 17916 5468
rect 17852 5408 17916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 10732 5068 10796 5132
rect 11952 4924 12016 4928
rect 11952 4868 11956 4924
rect 11956 4868 12012 4924
rect 12012 4868 12016 4924
rect 11952 4864 12016 4868
rect 12032 4924 12096 4928
rect 12032 4868 12036 4924
rect 12036 4868 12092 4924
rect 12092 4868 12096 4924
rect 12032 4864 12096 4868
rect 12112 4924 12176 4928
rect 12112 4868 12116 4924
rect 12116 4868 12172 4924
rect 12172 4868 12176 4924
rect 12112 4864 12176 4868
rect 12192 4924 12256 4928
rect 12192 4868 12196 4924
rect 12196 4868 12252 4924
rect 12252 4868 12256 4924
rect 12192 4864 12256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 11284 4796 11348 4860
rect 6684 4660 6748 4724
rect 2452 4524 2516 4588
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 17612 4380 17676 4384
rect 17612 4324 17616 4380
rect 17616 4324 17672 4380
rect 17672 4324 17676 4380
rect 17612 4320 17676 4324
rect 17692 4380 17756 4384
rect 17692 4324 17696 4380
rect 17696 4324 17752 4380
rect 17752 4324 17756 4380
rect 17692 4320 17756 4324
rect 17772 4380 17836 4384
rect 17772 4324 17776 4380
rect 17776 4324 17832 4380
rect 17832 4324 17836 4380
rect 17772 4320 17836 4324
rect 17852 4380 17916 4384
rect 17852 4324 17856 4380
rect 17856 4324 17912 4380
rect 17912 4324 17916 4380
rect 17852 4320 17916 4324
rect 9812 4252 9876 4316
rect 5948 3980 6012 4044
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 11952 3836 12016 3840
rect 11952 3780 11956 3836
rect 11956 3780 12012 3836
rect 12012 3780 12016 3836
rect 11952 3776 12016 3780
rect 12032 3836 12096 3840
rect 12032 3780 12036 3836
rect 12036 3780 12092 3836
rect 12092 3780 12096 3836
rect 12032 3776 12096 3780
rect 12112 3836 12176 3840
rect 12112 3780 12116 3836
rect 12116 3780 12172 3836
rect 12172 3780 12176 3836
rect 12112 3776 12176 3780
rect 12192 3836 12256 3840
rect 12192 3780 12196 3836
rect 12196 3780 12252 3836
rect 12252 3780 12256 3836
rect 12192 3776 12256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 4660 3572 4724 3636
rect 5396 3436 5460 3500
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 17612 3292 17676 3296
rect 17612 3236 17616 3292
rect 17616 3236 17672 3292
rect 17672 3236 17676 3292
rect 17612 3232 17676 3236
rect 17692 3292 17756 3296
rect 17692 3236 17696 3292
rect 17696 3236 17752 3292
rect 17752 3236 17756 3292
rect 17692 3232 17756 3236
rect 17772 3292 17836 3296
rect 17772 3236 17776 3292
rect 17776 3236 17832 3292
rect 17832 3236 17836 3292
rect 17772 3232 17836 3236
rect 17852 3292 17916 3296
rect 17852 3236 17856 3292
rect 17856 3236 17912 3292
rect 17912 3236 17916 3292
rect 17852 3232 17916 3236
rect 10916 3224 10980 3228
rect 10916 3168 10966 3224
rect 10966 3168 10980 3224
rect 10916 3164 10980 3168
rect 16620 2892 16684 2956
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 11952 2748 12016 2752
rect 11952 2692 11956 2748
rect 11956 2692 12012 2748
rect 12012 2692 12016 2748
rect 11952 2688 12016 2692
rect 12032 2748 12096 2752
rect 12032 2692 12036 2748
rect 12036 2692 12092 2748
rect 12092 2692 12096 2748
rect 12032 2688 12096 2692
rect 12112 2748 12176 2752
rect 12112 2692 12116 2748
rect 12116 2692 12172 2748
rect 12172 2692 12176 2748
rect 12112 2688 12176 2692
rect 12192 2748 12256 2752
rect 12192 2692 12196 2748
rect 12196 2692 12252 2748
rect 12252 2692 12256 2748
rect 12192 2688 12256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 9260 2620 9324 2684
rect 15884 2484 15948 2548
rect 6500 2348 6564 2412
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 17612 2204 17676 2208
rect 17612 2148 17616 2204
rect 17616 2148 17672 2204
rect 17672 2148 17676 2204
rect 17612 2144 17676 2148
rect 17692 2204 17756 2208
rect 17692 2148 17696 2204
rect 17696 2148 17752 2204
rect 17752 2148 17756 2204
rect 17692 2144 17756 2148
rect 17772 2204 17836 2208
rect 17772 2148 17776 2204
rect 17776 2148 17832 2204
rect 17832 2148 17836 2204
rect 17772 2144 17836 2148
rect 17852 2204 17916 2208
rect 17852 2148 17856 2204
rect 17856 2148 17912 2204
rect 17912 2148 17916 2204
rect 17852 2144 17916 2148
<< metal4 >>
rect 1944 16896 2264 17456
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 13294 2264 13568
rect 1944 13058 1986 13294
rect 2222 13058 2264 13294
rect 1944 12544 2264 13058
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 2604 17440 2924 17456
rect 2604 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2924 17440
rect 2604 16352 2924 17376
rect 5947 17100 6013 17101
rect 5947 17036 5948 17100
rect 6012 17036 6013 17100
rect 5947 17035 6013 17036
rect 2604 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2924 16352
rect 2604 15264 2924 16288
rect 4659 16012 4725 16013
rect 4659 15948 4660 16012
rect 4724 15948 4725 16012
rect 4659 15947 4725 15948
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2604 14176 2924 15200
rect 3923 14380 3989 14381
rect 3923 14316 3924 14380
rect 3988 14316 3989 14380
rect 3923 14315 3989 14316
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13954 2924 14112
rect 2604 13718 2646 13954
rect 2882 13718 2924 13954
rect 2604 13088 2924 13718
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2604 10912 2924 11936
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 3926 10845 3986 14315
rect 3923 10844 3989 10845
rect 3923 10780 3924 10844
rect 3988 10780 3989 10844
rect 3923 10779 3989 10780
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2451 8940 2517 8941
rect 2451 8876 2452 8940
rect 2516 8876 2517 8940
rect 2451 8875 2517 8876
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 2454 4589 2514 8875
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 3926 7853 3986 10779
rect 3923 7852 3989 7853
rect 3923 7788 3924 7852
rect 3988 7788 3989 7852
rect 3923 7787 3989 7788
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2451 4588 2517 4589
rect 2451 4524 2452 4588
rect 2516 4524 2517 4588
rect 2451 4523 2517 4524
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 4662 3637 4722 15947
rect 5395 12748 5461 12749
rect 5395 12684 5396 12748
rect 5460 12684 5461 12748
rect 5395 12683 5461 12684
rect 4659 3636 4725 3637
rect 4659 3572 4660 3636
rect 4724 3572 4725 3636
rect 4659 3571 4725 3572
rect 5398 3501 5458 12683
rect 5950 4045 6010 17035
rect 6944 16896 7264 17456
rect 6944 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7264 16896
rect 6944 15808 7264 16832
rect 6944 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7264 15808
rect 6499 15468 6565 15469
rect 6499 15404 6500 15468
rect 6564 15404 6565 15468
rect 6499 15403 6565 15404
rect 6131 13836 6197 13837
rect 6131 13772 6132 13836
rect 6196 13772 6197 13836
rect 6131 13771 6197 13772
rect 6134 6901 6194 13771
rect 6131 6900 6197 6901
rect 6131 6836 6132 6900
rect 6196 6836 6197 6900
rect 6131 6835 6197 6836
rect 5947 4044 6013 4045
rect 5947 3980 5948 4044
rect 6012 3980 6013 4044
rect 5947 3979 6013 3980
rect 5395 3500 5461 3501
rect 5395 3436 5396 3500
rect 5460 3436 5461 3500
rect 5395 3435 5461 3436
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 6502 2413 6562 15403
rect 6683 15332 6749 15333
rect 6683 15268 6684 15332
rect 6748 15268 6749 15332
rect 6683 15267 6749 15268
rect 6686 4725 6746 15267
rect 6944 14720 7264 15744
rect 6944 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7264 14720
rect 6944 13632 7264 14656
rect 6944 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7264 13632
rect 6944 13294 7264 13568
rect 6944 13058 6986 13294
rect 7222 13058 7264 13294
rect 7604 17440 7924 17456
rect 7604 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7924 17440
rect 7604 16352 7924 17376
rect 11944 16896 12264 17456
rect 11944 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12264 16896
rect 11099 16692 11165 16693
rect 11099 16628 11100 16692
rect 11164 16628 11165 16692
rect 11099 16627 11165 16628
rect 7604 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7924 16352
rect 7604 15264 7924 16288
rect 9259 15604 9325 15605
rect 9259 15540 9260 15604
rect 9324 15540 9325 15604
rect 9259 15539 9325 15540
rect 7604 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7924 15264
rect 7604 14176 7924 15200
rect 7604 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7924 14176
rect 7604 13954 7924 14112
rect 7604 13718 7646 13954
rect 7882 13718 7924 13954
rect 8155 13972 8221 13973
rect 8155 13908 8156 13972
rect 8220 13908 8221 13972
rect 8155 13907 8221 13908
rect 7419 13292 7485 13293
rect 7419 13228 7420 13292
rect 7484 13228 7485 13292
rect 7419 13227 7485 13228
rect 6944 12544 7264 13058
rect 6944 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7264 12544
rect 6944 11456 7264 12480
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 6944 10368 7264 11392
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6944 9280 7264 10304
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 7422 8397 7482 13227
rect 7604 13088 7924 13718
rect 7604 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7924 13088
rect 7604 12000 7924 13024
rect 8158 12341 8218 13907
rect 9075 13564 9141 13565
rect 9075 13500 9076 13564
rect 9140 13500 9141 13564
rect 9075 13499 9141 13500
rect 8155 12340 8221 12341
rect 8155 12276 8156 12340
rect 8220 12276 8221 12340
rect 8155 12275 8221 12276
rect 7604 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7924 12000
rect 7604 10912 7924 11936
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7604 9824 7924 10848
rect 9078 10301 9138 13499
rect 9262 13157 9322 15539
rect 9443 15332 9509 15333
rect 9443 15268 9444 15332
rect 9508 15268 9509 15332
rect 9443 15267 9509 15268
rect 10363 15332 10429 15333
rect 10363 15268 10364 15332
rect 10428 15268 10429 15332
rect 10363 15267 10429 15268
rect 10731 15332 10797 15333
rect 10731 15268 10732 15332
rect 10796 15268 10797 15332
rect 10731 15267 10797 15268
rect 10915 15332 10981 15333
rect 10915 15268 10916 15332
rect 10980 15268 10981 15332
rect 10915 15267 10981 15268
rect 9259 13156 9325 13157
rect 9259 13092 9260 13156
rect 9324 13092 9325 13156
rect 9259 13091 9325 13092
rect 9075 10300 9141 10301
rect 9075 10236 9076 10300
rect 9140 10236 9141 10300
rect 9075 10235 9141 10236
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7419 8396 7485 8397
rect 7419 8332 7420 8396
rect 7484 8332 7485 8396
rect 7419 8331 7485 8332
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 6944 7104 7264 8058
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 6683 4724 6749 4725
rect 6683 4660 6684 4724
rect 6748 4660 6749 4724
rect 6683 4659 6749 4660
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6499 2412 6565 2413
rect 6499 2348 6500 2412
rect 6564 2348 6565 2412
rect 6499 2347 6565 2348
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 2128 7264 2688
rect 7604 7648 7924 8672
rect 8155 7852 8221 7853
rect 8155 7788 8156 7852
rect 8220 7788 8221 7852
rect 8155 7787 8221 7788
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 8158 6357 8218 7787
rect 8155 6356 8221 6357
rect 8155 6292 8156 6356
rect 8220 6292 8221 6356
rect 8155 6291 8221 6292
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 9262 2685 9322 13091
rect 9446 5813 9506 15267
rect 9811 14788 9877 14789
rect 9811 14724 9812 14788
rect 9876 14724 9877 14788
rect 9811 14723 9877 14724
rect 9814 14650 9874 14723
rect 9814 14590 10058 14650
rect 9998 14517 10058 14590
rect 9995 14516 10061 14517
rect 9995 14452 9996 14516
rect 10060 14452 10061 14516
rect 9995 14451 10061 14452
rect 10366 11933 10426 15267
rect 10547 14788 10613 14789
rect 10547 14724 10548 14788
rect 10612 14724 10613 14788
rect 10547 14723 10613 14724
rect 10363 11932 10429 11933
rect 10363 11868 10364 11932
rect 10428 11868 10429 11932
rect 10363 11867 10429 11868
rect 9627 10300 9693 10301
rect 9627 10236 9628 10300
rect 9692 10236 9693 10300
rect 9627 10235 9693 10236
rect 9630 9690 9690 10235
rect 10550 9893 10610 14723
rect 10547 9892 10613 9893
rect 10547 9828 10548 9892
rect 10612 9828 10613 9892
rect 10547 9827 10613 9828
rect 9630 9630 9874 9690
rect 9814 7309 9874 9630
rect 9811 7308 9877 7309
rect 9811 7244 9812 7308
rect 9876 7244 9877 7308
rect 9811 7243 9877 7244
rect 9443 5812 9509 5813
rect 9443 5748 9444 5812
rect 9508 5748 9509 5812
rect 9443 5747 9509 5748
rect 9814 4317 9874 7243
rect 10734 5133 10794 15267
rect 10731 5132 10797 5133
rect 10731 5068 10732 5132
rect 10796 5068 10797 5132
rect 10731 5067 10797 5068
rect 9811 4316 9877 4317
rect 9811 4252 9812 4316
rect 9876 4252 9877 4316
rect 9811 4251 9877 4252
rect 10918 3229 10978 15267
rect 11102 12450 11162 16627
rect 11944 15808 12264 16832
rect 11944 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12264 15808
rect 11944 14720 12264 15744
rect 11944 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12264 14720
rect 11944 13632 12264 14656
rect 11944 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12264 13632
rect 11944 13294 12264 13568
rect 11944 13058 11986 13294
rect 12222 13058 12264 13294
rect 11944 12544 12264 13058
rect 11944 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12264 12544
rect 11102 12390 11346 12450
rect 11099 11388 11165 11389
rect 11099 11324 11100 11388
rect 11164 11324 11165 11388
rect 11099 11323 11165 11324
rect 11102 5677 11162 11323
rect 11099 5676 11165 5677
rect 11099 5612 11100 5676
rect 11164 5612 11165 5676
rect 11099 5611 11165 5612
rect 11286 4861 11346 12390
rect 11651 11932 11717 11933
rect 11651 11868 11652 11932
rect 11716 11868 11717 11932
rect 11651 11867 11717 11868
rect 11654 10845 11714 11867
rect 11944 11456 12264 12480
rect 11944 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12264 11456
rect 11651 10844 11717 10845
rect 11651 10780 11652 10844
rect 11716 10780 11717 10844
rect 11651 10779 11717 10780
rect 11944 10368 12264 11392
rect 11944 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12264 10368
rect 11944 9280 12264 10304
rect 12604 17440 12924 17456
rect 12604 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12924 17440
rect 12604 16352 12924 17376
rect 16944 16896 17264 17456
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 14411 16420 14477 16421
rect 14411 16356 14412 16420
rect 14476 16356 14477 16420
rect 14411 16355 14477 16356
rect 12604 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12924 16352
rect 12604 15264 12924 16288
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12604 14176 12924 15200
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12604 13954 12924 14112
rect 12604 13718 12646 13954
rect 12882 13718 12924 13954
rect 13491 13836 13557 13837
rect 13491 13772 13492 13836
rect 13556 13772 13557 13836
rect 13491 13771 13557 13772
rect 12604 13088 12924 13718
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12604 12000 12924 13024
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12387 10300 12453 10301
rect 12387 10236 12388 10300
rect 12452 10236 12453 10300
rect 12387 10235 12453 10236
rect 12390 9893 12450 10235
rect 12387 9892 12453 9893
rect 12387 9828 12388 9892
rect 12452 9828 12453 9892
rect 12387 9827 12453 9828
rect 11944 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12264 9280
rect 11944 8294 12264 9216
rect 11944 8192 11986 8294
rect 12222 8192 12264 8294
rect 11944 8128 11952 8192
rect 12256 8128 12264 8192
rect 11944 8058 11986 8128
rect 12222 8058 12264 8128
rect 11944 7104 12264 8058
rect 11944 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12264 7104
rect 11944 6016 12264 7040
rect 11944 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12264 6016
rect 11944 4928 12264 5952
rect 11944 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12264 4928
rect 11283 4860 11349 4861
rect 11283 4796 11284 4860
rect 11348 4796 11349 4860
rect 11283 4795 11349 4796
rect 11944 3840 12264 4864
rect 11944 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12264 3840
rect 11944 3294 12264 3776
rect 10915 3228 10981 3229
rect 10915 3164 10916 3228
rect 10980 3164 10981 3228
rect 10915 3163 10981 3164
rect 11944 3058 11986 3294
rect 12222 3058 12264 3294
rect 11944 2752 12264 3058
rect 11944 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12264 2752
rect 9259 2684 9325 2685
rect 9259 2620 9260 2684
rect 9324 2620 9325 2684
rect 9259 2619 9325 2620
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
rect 11944 2128 12264 2688
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12604 8954 12924 9760
rect 12604 8736 12646 8954
rect 12882 8736 12924 8954
rect 12604 8672 12612 8736
rect 12676 8672 12692 8718
rect 12756 8672 12772 8718
rect 12836 8672 12852 8718
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 13494 8533 13554 13771
rect 13675 13428 13741 13429
rect 13675 13364 13676 13428
rect 13740 13364 13741 13428
rect 13675 13363 13741 13364
rect 13491 8532 13557 8533
rect 13491 8468 13492 8532
rect 13556 8468 13557 8532
rect 13491 8467 13557 8468
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12604 6560 12924 7584
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12604 5472 12924 6496
rect 13678 6493 13738 13363
rect 14414 6901 14474 16355
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16619 15604 16685 15605
rect 16619 15540 16620 15604
rect 16684 15540 16685 15604
rect 16619 15539 16685 15540
rect 15331 14380 15397 14381
rect 15331 14316 15332 14380
rect 15396 14316 15397 14380
rect 15331 14315 15397 14316
rect 14963 13836 15029 13837
rect 14963 13772 14964 13836
rect 15028 13772 15029 13836
rect 14963 13771 15029 13772
rect 14966 8941 15026 13771
rect 15147 10980 15213 10981
rect 15147 10916 15148 10980
rect 15212 10916 15213 10980
rect 15147 10915 15213 10916
rect 14963 8940 15029 8941
rect 14963 8876 14964 8940
rect 15028 8876 15029 8940
rect 14963 8875 15029 8876
rect 14411 6900 14477 6901
rect 14411 6836 14412 6900
rect 14476 6836 14477 6900
rect 14411 6835 14477 6836
rect 13675 6492 13741 6493
rect 13675 6428 13676 6492
rect 13740 6428 13741 6492
rect 13675 6427 13741 6428
rect 14966 6221 15026 8875
rect 15150 6901 15210 10915
rect 15334 8261 15394 14315
rect 15883 13564 15949 13565
rect 15883 13500 15884 13564
rect 15948 13500 15949 13564
rect 15883 13499 15949 13500
rect 15331 8260 15397 8261
rect 15331 8196 15332 8260
rect 15396 8196 15397 8260
rect 15331 8195 15397 8196
rect 15147 6900 15213 6901
rect 15147 6836 15148 6900
rect 15212 6836 15213 6900
rect 15147 6835 15213 6836
rect 14963 6220 15029 6221
rect 14963 6156 14964 6220
rect 15028 6156 15029 6220
rect 14963 6155 15029 6156
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12604 4384 12924 5408
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3954 12924 4320
rect 12604 3718 12646 3954
rect 12882 3718 12924 3954
rect 12604 3296 12924 3718
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 15886 2549 15946 13499
rect 16622 2957 16682 15539
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13294 17264 13568
rect 16944 13058 16986 13294
rect 17222 13058 17264 13294
rect 16803 12748 16869 12749
rect 16803 12684 16804 12748
rect 16868 12684 16869 12748
rect 16803 12683 16869 12684
rect 16806 10029 16866 12683
rect 16944 12544 17264 13058
rect 17604 17440 17924 17456
rect 17604 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17924 17440
rect 17604 16352 17924 17376
rect 17604 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17924 16352
rect 17604 15264 17924 16288
rect 17604 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17924 15264
rect 17604 14176 17924 15200
rect 17604 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17924 14176
rect 17604 13954 17924 14112
rect 17604 13718 17646 13954
rect 17882 13718 17924 13954
rect 17604 13088 17924 13718
rect 17604 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17924 13088
rect 17355 12748 17421 12749
rect 17355 12684 17356 12748
rect 17420 12684 17421 12748
rect 17355 12683 17421 12684
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 17358 12341 17418 12683
rect 17355 12340 17421 12341
rect 17355 12276 17356 12340
rect 17420 12276 17421 12340
rect 17355 12275 17421 12276
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16803 10028 16869 10029
rect 16803 9964 16804 10028
rect 16868 9964 16869 10028
rect 16803 9963 16869 9964
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8294 17264 9216
rect 16944 8192 16986 8294
rect 17222 8192 17264 8294
rect 16944 8128 16952 8192
rect 17256 8128 17264 8192
rect 16944 8058 16986 8128
rect 17222 8058 17264 8128
rect 16944 7104 17264 8058
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3294 17264 3776
rect 16944 3058 16986 3294
rect 17222 3058 17264 3294
rect 16619 2956 16685 2957
rect 16619 2892 16620 2956
rect 16684 2892 16685 2956
rect 16619 2891 16685 2892
rect 16944 2752 17264 3058
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 15883 2548 15949 2549
rect 15883 2484 15884 2548
rect 15948 2484 15949 2548
rect 15883 2483 15949 2484
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 16944 2128 17264 2688
rect 17604 12000 17924 13024
rect 17604 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17924 12000
rect 17604 10912 17924 11936
rect 17604 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17924 10912
rect 17604 9824 17924 10848
rect 17604 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17924 9824
rect 17604 8954 17924 9760
rect 17604 8736 17646 8954
rect 17882 8736 17924 8954
rect 17604 8672 17612 8736
rect 17676 8672 17692 8718
rect 17756 8672 17772 8718
rect 17836 8672 17852 8718
rect 17916 8672 17924 8736
rect 17604 7648 17924 8672
rect 17604 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17924 7648
rect 17604 6560 17924 7584
rect 17604 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17924 6560
rect 17604 5472 17924 6496
rect 17604 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17924 5472
rect 17604 4384 17924 5408
rect 17604 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17924 4384
rect 17604 3954 17924 4320
rect 17604 3718 17646 3954
rect 17882 3718 17924 3954
rect 17604 3296 17924 3718
rect 17604 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17924 3296
rect 17604 2208 17924 3232
rect 17604 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17924 2208
rect 17604 2128 17924 2144
<< via4 >>
rect 1986 13058 2222 13294
rect 2646 13718 2882 13954
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 1986 3058 2222 3294
rect 2646 3718 2882 3954
rect 6986 13058 7222 13294
rect 7646 13718 7882 13954
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 6986 3058 7222 3294
rect 7646 3718 7882 3954
rect 11986 13058 12222 13294
rect 12646 13718 12882 13954
rect 11986 8192 12222 8294
rect 11986 8128 12016 8192
rect 12016 8128 12032 8192
rect 12032 8128 12096 8192
rect 12096 8128 12112 8192
rect 12112 8128 12176 8192
rect 12176 8128 12192 8192
rect 12192 8128 12222 8192
rect 11986 8058 12222 8128
rect 11986 3058 12222 3294
rect 12646 8736 12882 8954
rect 12646 8718 12676 8736
rect 12676 8718 12692 8736
rect 12692 8718 12756 8736
rect 12756 8718 12772 8736
rect 12772 8718 12836 8736
rect 12836 8718 12852 8736
rect 12852 8718 12882 8736
rect 12646 3718 12882 3954
rect 16986 13058 17222 13294
rect 17646 13718 17882 13954
rect 16986 8192 17222 8294
rect 16986 8128 17016 8192
rect 17016 8128 17032 8192
rect 17032 8128 17096 8192
rect 17096 8128 17112 8192
rect 17112 8128 17176 8192
rect 17176 8128 17192 8192
rect 17192 8128 17222 8192
rect 16986 8058 17222 8128
rect 16986 3058 17222 3294
rect 17646 8736 17882 8954
rect 17646 8718 17676 8736
rect 17676 8718 17692 8736
rect 17692 8718 17756 8736
rect 17756 8718 17772 8736
rect 17772 8718 17836 8736
rect 17836 8718 17852 8736
rect 17852 8718 17882 8736
rect 17646 3718 17882 3954
<< metal5 >>
rect 1056 13954 18908 13996
rect 1056 13718 2646 13954
rect 2882 13718 7646 13954
rect 7882 13718 12646 13954
rect 12882 13718 17646 13954
rect 17882 13718 18908 13954
rect 1056 13676 18908 13718
rect 1056 13294 18908 13336
rect 1056 13058 1986 13294
rect 2222 13058 6986 13294
rect 7222 13058 11986 13294
rect 12222 13058 16986 13294
rect 17222 13058 18908 13294
rect 1056 13016 18908 13058
rect 1056 8954 18908 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 12646 8954
rect 12882 8718 17646 8954
rect 17882 8718 18908 8954
rect 1056 8676 18908 8718
rect 1056 8294 18908 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 11986 8294
rect 12222 8058 16986 8294
rect 17222 8058 18908 8294
rect 1056 8016 18908 8058
rect 1056 3954 18908 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 12646 3954
rect 12882 3718 17646 3954
rect 17882 3718 18908 3954
rect 1056 3676 18908 3718
rect 1056 3294 18908 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 11986 3294
rect 12222 3058 16986 3294
rect 17222 3058 18908 3294
rect 1056 3016 18908 3058
use sky130_fd_sc_hd__inv_2  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16928 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17296 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13524 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11868 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9384 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _175_
timestamp 1704896540
transform 1 0 2116 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _177_
timestamp 1704896540
transform 1 0 11408 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _178_
timestamp 1704896540
transform 1 0 2116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _179_
timestamp 1704896540
transform -1 0 13340 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _180_
timestamp 1704896540
transform 1 0 2484 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4140 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17572 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _183_
timestamp 1704896540
transform 1 0 12604 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _184_
timestamp 1704896540
transform -1 0 5520 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_4  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16836 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9844 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_4  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14720 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__xnor2_4  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12052 0 1 4352
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _189_
timestamp 1704896540
transform 1 0 2392 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18216 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _191_
timestamp 1704896540
transform 1 0 15088 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7820 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _194_
timestamp 1704896540
transform 1 0 2944 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _195_
timestamp 1704896540
transform 1 0 2576 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10396 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16652 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18400 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _199_
timestamp 1704896540
transform -1 0 13248 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13892 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp 1704896540
transform 1 0 4968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15272 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15548 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_1  _205_
timestamp 1704896540
transform -1 0 15088 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11408 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _207_
timestamp 1704896540
transform 1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _208_
timestamp 1704896540
transform -1 0 13800 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _209_
timestamp 1704896540
transform 1 0 12512 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_1  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16468 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _211_
timestamp 1704896540
transform 1 0 4784 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _212_
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _213_
timestamp 1704896540
transform 1 0 5152 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _214_
timestamp 1704896540
transform 1 0 3128 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _215_
timestamp 1704896540
transform 1 0 4968 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_1  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _217_
timestamp 1704896540
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15272 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _220_
timestamp 1704896540
transform -1 0 13616 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _222_
timestamp 1704896540
transform 1 0 5428 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _223_
timestamp 1704896540
transform 1 0 17756 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12236 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _225_
timestamp 1704896540
transform -1 0 3312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _226_
timestamp 1704896540
transform -1 0 14996 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _227_
timestamp 1704896540
transform 1 0 16652 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10672 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9752 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _230_
timestamp 1704896540
transform -1 0 7820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _231_
timestamp 1704896540
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2668 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16744 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10120 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_4  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13248 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__o31a_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _237_
timestamp 1704896540
transform 1 0 14536 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _238_
timestamp 1704896540
transform -1 0 8372 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14720 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _240_
timestamp 1704896540
transform -1 0 9660 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _241_
timestamp 1704896540
transform 1 0 4232 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _242_
timestamp 1704896540
transform 1 0 4048 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _243_
timestamp 1704896540
transform -1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12420 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2668 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _246_
timestamp 1704896540
transform -1 0 10212 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7084 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _248_
timestamp 1704896540
transform -1 0 4600 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _249_
timestamp 1704896540
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _250_
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _252_
timestamp 1704896540
transform -1 0 7268 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _253_
timestamp 1704896540
transform -1 0 4140 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _254_
timestamp 1704896540
transform 1 0 17940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _255_
timestamp 1704896540
transform 1 0 15732 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _256_
timestamp 1704896540
transform -1 0 9200 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_4  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14536 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__a21o_1  _258_
timestamp 1704896540
transform -1 0 8740 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16468 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _260_
timestamp 1704896540
transform -1 0 12696 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _261_
timestamp 1704896540
transform -1 0 14720 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _262_
timestamp 1704896540
transform -1 0 13616 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _263_
timestamp 1704896540
transform -1 0 14628 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _264_
timestamp 1704896540
transform 1 0 15916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _266_
timestamp 1704896540
transform -1 0 18124 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17112 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7452 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _269_
timestamp 1704896540
transform -1 0 10580 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5520 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _271_
timestamp 1704896540
transform 1 0 12420 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _272_
timestamp 1704896540
transform -1 0 3588 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1704896540
transform -1 0 7084 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _274_
timestamp 1704896540
transform -1 0 14720 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _275_
timestamp 1704896540
transform 1 0 15180 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_4  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4968 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _277_
timestamp 1704896540
transform 1 0 9108 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _278_
timestamp 1704896540
transform -1 0 17388 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _279_
timestamp 1704896540
transform 1 0 3772 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _280_
timestamp 1704896540
transform -1 0 2576 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp 1704896540
transform 1 0 8096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _282_
timestamp 1704896540
transform -1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _283_
timestamp 1704896540
transform -1 0 3680 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _284_
timestamp 1704896540
transform -1 0 7360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _285_
timestamp 1704896540
transform 1 0 8096 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _286_
timestamp 1704896540
transform 1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _287_
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _288_
timestamp 1704896540
transform 1 0 3404 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7636 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _290_
timestamp 1704896540
transform -1 0 6256 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _291_
timestamp 1704896540
transform -1 0 16652 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _292_
timestamp 1704896540
transform -1 0 12696 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _293_
timestamp 1704896540
transform -1 0 15088 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _294_
timestamp 1704896540
transform -1 0 8648 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _295_
timestamp 1704896540
transform -1 0 18584 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _296_
timestamp 1704896540
transform 1 0 5888 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _297_
timestamp 1704896540
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _298_
timestamp 1704896540
transform -1 0 14628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7728 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14628 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _302_
timestamp 1704896540
transform -1 0 18032 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _303_
timestamp 1704896540
transform -1 0 15548 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _304_
timestamp 1704896540
transform 1 0 17940 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _305_
timestamp 1704896540
transform 1 0 13432 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _306_
timestamp 1704896540
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _307_
timestamp 1704896540
transform -1 0 9292 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _308_
timestamp 1704896540
transform 1 0 1472 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _309_
timestamp 1704896540
transform -1 0 14444 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _310_
timestamp 1704896540
transform 1 0 9660 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14720 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _312_
timestamp 1704896540
transform -1 0 9936 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _313_
timestamp 1704896540
transform -1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _314_
timestamp 1704896540
transform -1 0 16376 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _315_
timestamp 1704896540
transform -1 0 5888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _316_
timestamp 1704896540
transform 1 0 14076 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _319_
timestamp 1704896540
transform 1 0 15640 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _320_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14352 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _321_
timestamp 1704896540
transform -1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _322_
timestamp 1704896540
transform -1 0 8648 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _323_
timestamp 1704896540
transform 1 0 16744 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _324_
timestamp 1704896540
transform 1 0 7728 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_2  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2392 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _326_
timestamp 1704896540
transform -1 0 15364 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _327_
timestamp 1704896540
transform 1 0 9936 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _328_
timestamp 1704896540
transform -1 0 15272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _329_
timestamp 1704896540
transform 1 0 10396 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10396 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _331_
timestamp 1704896540
transform 1 0 1472 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _332_
timestamp 1704896540
transform 1 0 16652 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _333_
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _334_
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11960 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _336_
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _337_
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _338_
timestamp 1704896540
transform -1 0 14812 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _339_
timestamp 1704896540
transform -1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _340_
timestamp 1704896540
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _341_
timestamp 1704896540
transform -1 0 7176 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _342_
timestamp 1704896540
transform -1 0 7728 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _343_
timestamp 1704896540
transform 1 0 13156 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _344_
timestamp 1704896540
transform -1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _345_
timestamp 1704896540
transform 1 0 14076 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _346_
timestamp 1704896540
transform -1 0 7360 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _347_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15088 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1704896540
transform 1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__nand3b_2  clone1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2392 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26
timestamp 1704896540
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_35
timestamp 1704896540
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_88
timestamp 1704896540
transform 1 0 9200 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_96
timestamp 1704896540
transform 1 0 9936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_103
timestamp 1704896540
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1704896540
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15180 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_164 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_173
timestamp 1704896540
transform 1 0 17020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_179
timestamp 1704896540
transform 1 0 17572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_185
timestamp 1704896540
transform 1 0 18124 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_14
timestamp 1704896540
transform 1 0 2392 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_26
timestamp 1704896540
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_33
timestamp 1704896540
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_45
timestamp 1704896540
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_53
timestamp 1704896540
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_90
timestamp 1704896540
transform 1 0 9384 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_102
timestamp 1704896540
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_117
timestamp 1704896540
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_126
timestamp 1704896540
transform 1 0 12696 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_138
timestamp 1704896540
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_142
timestamp 1704896540
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_147
timestamp 1704896540
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_159
timestamp 1704896540
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_189
timestamp 1704896540
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_36
timestamp 1704896540
transform 1 0 4416 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_48
timestamp 1704896540
transform 1 0 5520 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_60
timestamp 1704896540
transform 1 0 6624 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_72
timestamp 1704896540
transform 1 0 7728 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_91
timestamp 1704896540
transform 1 0 9476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_103
timestamp 1704896540
transform 1 0 10580 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_115
timestamp 1704896540
transform 1 0 11684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_127
timestamp 1704896540
transform 1 0 12788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_141
timestamp 1704896540
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_155
timestamp 1704896540
transform 1 0 15364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_167
timestamp 1704896540
transform 1 0 16468 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_179
timestamp 1704896540
transform 1 0 17572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_187
timestamp 1704896540
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_7
timestamp 1704896540
transform 1 0 1748 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_24
timestamp 1704896540
transform 1 0 3312 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_36
timestamp 1704896540
transform 1 0 4416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_48
timestamp 1704896540
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 1704896540
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_102
timestamp 1704896540
transform 1 0 10488 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1704896540
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13708 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_143
timestamp 1704896540
transform 1 0 14260 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_175
timestamp 1704896540
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_181
timestamp 1704896540
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_185
timestamp 1704896540
transform 1 0 18124 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1704896540
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_92
timestamp 1704896540
transform 1 0 9568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_96
timestamp 1704896540
transform 1 0 9936 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_125
timestamp 1704896540
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_137
timestamp 1704896540
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_148
timestamp 1704896540
transform 1 0 14720 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_156
timestamp 1704896540
transform 1 0 15456 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_160
timestamp 1704896540
transform 1 0 15824 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_173
timestamp 1704896540
transform 1 0 17020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_185
timestamp 1704896540
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_189
timestamp 1704896540
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_7
timestamp 1704896540
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_17
timestamp 1704896540
transform 1 0 2668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_29
timestamp 1704896540
transform 1 0 3772 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_37
timestamp 1704896540
transform 1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_46
timestamp 1704896540
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1704896540
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_69
timestamp 1704896540
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_77
timestamp 1704896540
transform 1 0 8188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_89
timestamp 1704896540
transform 1 0 9292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_101
timestamp 1704896540
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1704896540
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_123
timestamp 1704896540
transform 1 0 12420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_130
timestamp 1704896540
transform 1 0 13064 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_138
timestamp 1704896540
transform 1 0 13800 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_150
timestamp 1704896540
transform 1 0 14904 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_156
timestamp 1704896540
transform 1 0 15456 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_189
timestamp 1704896540
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_37
timestamp 1704896540
transform 1 0 4508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_49
timestamp 1704896540
transform 1 0 5612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_61
timestamp 1704896540
transform 1 0 6716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_73
timestamp 1704896540
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 1704896540
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_109
timestamp 1704896540
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_135
timestamp 1704896540
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_150
timestamp 1704896540
transform 1 0 14904 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_162
timestamp 1704896540
transform 1 0 16008 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_172
timestamp 1704896540
transform 1 0 16928 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_184
timestamp 1704896540
transform 1 0 18032 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_12
timestamp 1704896540
transform 1 0 2208 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_24
timestamp 1704896540
transform 1 0 3312 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_36
timestamp 1704896540
transform 1 0 4416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_48
timestamp 1704896540
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_65
timestamp 1704896540
transform 1 0 7084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_77
timestamp 1704896540
transform 1 0 8188 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_89
timestamp 1704896540
transform 1 0 9292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_95
timestamp 1704896540
transform 1 0 9844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_102
timestamp 1704896540
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1704896540
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_131
timestamp 1704896540
transform 1 0 13156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_138
timestamp 1704896540
transform 1 0 13800 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_150
timestamp 1704896540
transform 1 0 14904 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_158
timestamp 1704896540
transform 1 0 15640 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_181
timestamp 1704896540
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_185
timestamp 1704896540
transform 1 0 18124 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_23
timestamp 1704896540
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_45
timestamp 1704896540
transform 1 0 5244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_57
timestamp 1704896540
transform 1 0 6348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_69
timestamp 1704896540
transform 1 0 7452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1704896540
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_100
timestamp 1704896540
transform 1 0 10304 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_112
timestamp 1704896540
transform 1 0 11408 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_120
timestamp 1704896540
transform 1 0 12144 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_126
timestamp 1704896540
transform 1 0 12696 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1704896540
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_153
timestamp 1704896540
transform 1 0 15180 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_171
timestamp 1704896540
transform 1 0 16836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_183
timestamp 1704896540
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_7
timestamp 1704896540
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_19
timestamp 1704896540
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_31
timestamp 1704896540
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_43
timestamp 1704896540
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_69
timestamp 1704896540
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_80
timestamp 1704896540
transform 1 0 8464 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_92
timestamp 1704896540
transform 1 0 9568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_104
timestamp 1704896540
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_136
timestamp 1704896540
transform 1 0 13616 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_145
timestamp 1704896540
transform 1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_157
timestamp 1704896540
transform 1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1704896540
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_181
timestamp 1704896540
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_189
timestamp 1704896540
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_9
timestamp 1704896540
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_19
timestamp 1704896540
transform 1 0 2852 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_42
timestamp 1704896540
transform 1 0 4968 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_54
timestamp 1704896540
transform 1 0 6072 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_66
timestamp 1704896540
transform 1 0 7176 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_74
timestamp 1704896540
transform 1 0 7912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1704896540
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1704896540
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1704896540
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1704896540
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1704896540
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1704896540
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1704896540
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1704896540
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_177
timestamp 1704896540
transform 1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_183
timestamp 1704896540
transform 1 0 17940 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_189
timestamp 1704896540
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_13
timestamp 1704896540
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_32
timestamp 1704896540
transform 1 0 4048 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_38
timestamp 1704896540
transform 1 0 4600 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_50
timestamp 1704896540
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_71
timestamp 1704896540
transform 1 0 7636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_83
timestamp 1704896540
transform 1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_91
timestamp 1704896540
transform 1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_99
timestamp 1704896540
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1704896540
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_113
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_121
timestamp 1704896540
transform 1 0 12236 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1704896540
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_137
timestamp 1704896540
transform 1 0 13708 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_147
timestamp 1704896540
transform 1 0 14628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_159
timestamp 1704896540
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1704896540
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_181
timestamp 1704896540
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_189
timestamp 1704896540
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_12
timestamp 1704896540
transform 1 0 2208 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_24
timestamp 1704896540
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1704896540
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1704896540
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_88
timestamp 1704896540
transform 1 0 9200 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_100
timestamp 1704896540
transform 1 0 10304 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_112
timestamp 1704896540
transform 1 0 11408 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_124
timestamp 1704896540
transform 1 0 12512 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_136
timestamp 1704896540
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_141
timestamp 1704896540
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_157
timestamp 1704896540
transform 1 0 15548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_169
timestamp 1704896540
transform 1 0 16652 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_177
timestamp 1704896540
transform 1 0 17388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_6
timestamp 1704896540
transform 1 0 1656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_17
timestamp 1704896540
transform 1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_43
timestamp 1704896540
transform 1 0 5060 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1704896540
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1704896540
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1704896540
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1704896540
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1704896540
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1704896540
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1704896540
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1704896540
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_161
timestamp 1704896540
transform 1 0 15916 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_174
timestamp 1704896540
transform 1 0 17112 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_182
timestamp 1704896540
transform 1 0 17848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_189
timestamp 1704896540
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_7
timestamp 1704896540
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_11
timestamp 1704896540
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 1704896540
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_44
timestamp 1704896540
transform 1 0 5152 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_56
timestamp 1704896540
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_68
timestamp 1704896540
transform 1 0 7360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_80
timestamp 1704896540
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_97
timestamp 1704896540
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_108
timestamp 1704896540
transform 1 0 11040 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_117
timestamp 1704896540
transform 1 0 11868 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_129
timestamp 1704896540
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1704896540
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_141
timestamp 1704896540
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_158
timestamp 1704896540
transform 1 0 15640 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_187
timestamp 1704896540
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_8
timestamp 1704896540
transform 1 0 1840 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_46
timestamp 1704896540
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1704896540
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1704896540
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1704896540
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1704896540
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1704896540
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_144
timestamp 1704896540
transform 1 0 14352 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_156
timestamp 1704896540
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_181
timestamp 1704896540
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_185
timestamp 1704896540
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_7
timestamp 1704896540
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_17
timestamp 1704896540
transform 1 0 2668 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_25
timestamp 1704896540
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_33
timestamp 1704896540
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_47
timestamp 1704896540
transform 1 0 5428 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_51
timestamp 1704896540
transform 1 0 5796 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_57
timestamp 1704896540
transform 1 0 6348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_69
timestamp 1704896540
transform 1 0 7452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1704896540
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1704896540
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1704896540
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_125
timestamp 1704896540
transform 1 0 12604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1704896540
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_155
timestamp 1704896540
transform 1 0 15364 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1704896540
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1704896540
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_189
timestamp 1704896540
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_7
timestamp 1704896540
transform 1 0 1748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_19
timestamp 1704896540
transform 1 0 2852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_33
timestamp 1704896540
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_45
timestamp 1704896540
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1704896540
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_65
timestamp 1704896540
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_72
timestamp 1704896540
transform 1 0 7728 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_84
timestamp 1704896540
transform 1 0 8832 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_103
timestamp 1704896540
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1704896540
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_113
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_121
timestamp 1704896540
transform 1 0 12236 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_133
timestamp 1704896540
transform 1 0 13340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_141
timestamp 1704896540
transform 1 0 14076 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_148
timestamp 1704896540
transform 1 0 14720 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_160
timestamp 1704896540
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_184
timestamp 1704896540
transform 1 0 18032 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_17
timestamp 1704896540
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_25
timestamp 1704896540
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1704896540
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_68
timestamp 1704896540
transform 1 0 7360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_73
timestamp 1704896540
transform 1 0 7820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1704896540
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_89
timestamp 1704896540
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_94
timestamp 1704896540
transform 1 0 9752 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_105
timestamp 1704896540
transform 1 0 10764 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_111
timestamp 1704896540
transform 1 0 11316 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_121
timestamp 1704896540
transform 1 0 12236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1704896540
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_154
timestamp 1704896540
transform 1 0 15272 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_166
timestamp 1704896540
transform 1 0 16376 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_178
timestamp 1704896540
transform 1 0 17480 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_7
timestamp 1704896540
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_19
timestamp 1704896540
transform 1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1704896540
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_73
timestamp 1704896540
transform 1 0 7820 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_79
timestamp 1704896540
transform 1 0 8372 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_91
timestamp 1704896540
transform 1 0 9476 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_104
timestamp 1704896540
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_125
timestamp 1704896540
transform 1 0 12604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_133
timestamp 1704896540
transform 1 0 13340 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_141
timestamp 1704896540
transform 1 0 14076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_153
timestamp 1704896540
transform 1 0 15180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1704896540
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1704896540
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_181
timestamp 1704896540
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_189
timestamp 1704896540
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_15
timestamp 1704896540
transform 1 0 2484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_21
timestamp 1704896540
transform 1 0 3036 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1704896540
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_53
timestamp 1704896540
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_61
timestamp 1704896540
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1704896540
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1704896540
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1704896540
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_93
timestamp 1704896540
transform 1 0 9660 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_105
timestamp 1704896540
transform 1 0 10764 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_117
timestamp 1704896540
transform 1 0 11868 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_132
timestamp 1704896540
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_141
timestamp 1704896540
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_145
timestamp 1704896540
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_162
timestamp 1704896540
transform 1 0 16008 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_174
timestamp 1704896540
transform 1 0 17112 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_186
timestamp 1704896540
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_7
timestamp 1704896540
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_19
timestamp 1704896540
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_31
timestamp 1704896540
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_43
timestamp 1704896540
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1704896540
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_81
timestamp 1704896540
transform 1 0 8556 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_89
timestamp 1704896540
transform 1 0 9292 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_101
timestamp 1704896540
transform 1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 1704896540
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_126
timestamp 1704896540
transform 1 0 12696 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_134
timestamp 1704896540
transform 1 0 13432 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_140
timestamp 1704896540
transform 1 0 13984 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_152
timestamp 1704896540
transform 1 0 15088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_164
timestamp 1704896540
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_181
timestamp 1704896540
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_185
timestamp 1704896540
transform 1 0 18124 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1704896540
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1704896540
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1704896540
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1704896540
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1704896540
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1704896540
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_93
timestamp 1704896540
transform 1 0 9660 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_101
timestamp 1704896540
transform 1 0 10396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_113
timestamp 1704896540
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_125
timestamp 1704896540
transform 1 0 12604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1704896540
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 1704896540
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_145
timestamp 1704896540
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_159
timestamp 1704896540
transform 1 0 15732 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_167
timestamp 1704896540
transform 1 0 16468 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_175
timestamp 1704896540
transform 1 0 17204 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_187
timestamp 1704896540
transform 1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_7
timestamp 1704896540
transform 1 0 1748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_19
timestamp 1704896540
transform 1 0 2852 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1704896540
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4692 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_47
timestamp 1704896540
transform 1 0 5428 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_53
timestamp 1704896540
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1704896540
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_79
timestamp 1704896540
transform 1 0 8372 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_101
timestamp 1704896540
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1704896540
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1704896540
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_125
timestamp 1704896540
transform 1 0 12604 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_131
timestamp 1704896540
transform 1 0 13156 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_154
timestamp 1704896540
transform 1 0 15272 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1704896540
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_176
timestamp 1704896540
transform 1 0 17296 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_188
timestamp 1704896540
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1704896540
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1704896540
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_53
timestamp 1704896540
transform 1 0 5980 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_67
timestamp 1704896540
transform 1 0 7268 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_75
timestamp 1704896540
transform 1 0 8004 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 1704896540
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1704896540
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1704896540
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_97
timestamp 1704896540
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_108
timestamp 1704896540
transform 1 0 11040 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_120
timestamp 1704896540
transform 1 0 12144 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_148
timestamp 1704896540
transform 1 0 14720 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_157
timestamp 1704896540
transform 1 0 15548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_169
timestamp 1704896540
transform 1 0 16652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_177
timestamp 1704896540
transform 1 0 17388 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_189
timestamp 1704896540
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_3
timestamp 1704896540
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_12
timestamp 1704896540
transform 1 0 2208 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_36
timestamp 1704896540
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_48
timestamp 1704896540
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1704896540
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1704896540
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_81
timestamp 1704896540
transform 1 0 8556 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_96
timestamp 1704896540
transform 1 0 9936 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_108
timestamp 1704896540
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_113
timestamp 1704896540
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_123
timestamp 1704896540
transform 1 0 12420 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_136
timestamp 1704896540
transform 1 0 13616 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_148
timestamp 1704896540
transform 1 0 14720 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_160
timestamp 1704896540
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1704896540
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1704896540
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1704896540
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_35
timestamp 1704896540
transform 1 0 4324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_52
timestamp 1704896540
transform 1 0 5888 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_58
timestamp 1704896540
transform 1 0 6440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_66
timestamp 1704896540
transform 1 0 7176 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 1704896540
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_88
timestamp 1704896540
transform 1 0 9200 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_92
timestamp 1704896540
transform 1 0 9568 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_97
timestamp 1704896540
transform 1 0 10028 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_104
timestamp 1704896540
transform 1 0 10672 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_116
timestamp 1704896540
transform 1 0 11776 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1704896540
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_154
timestamp 1704896540
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_163
timestamp 1704896540
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_174
timestamp 1704896540
transform 1 0 17112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_178
timestamp 1704896540
transform 1 0 17480 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_188
timestamp 1704896540
transform 1 0 18400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_11
timestamp 1704896540
transform 1 0 2116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_20
timestamp 1704896540
transform 1 0 2944 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_29
timestamp 1704896540
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_41
timestamp 1704896540
transform 1 0 4876 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_48
timestamp 1704896540
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1704896540
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1704896540
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_81
timestamp 1704896540
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_85
timestamp 1704896540
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_97
timestamp 1704896540
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1704896540
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1704896540
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1704896540
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_137
timestamp 1704896540
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_141
timestamp 1704896540
transform 1 0 14076 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_147
timestamp 1704896540
transform 1 0 14628 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_163
timestamp 1704896540
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1704896540
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_181
timestamp 1704896540
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_185
timestamp 1704896540
transform 1 0 18124 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1704896540
transform 1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1704896540
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1704896540
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1704896540
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1704896540
transform 1 0 1840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1704896540
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1704896540
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1704896540
transform 1 0 18216 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1704896540
transform 1 0 17572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1704896540
transform 1 0 18216 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1704896540
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1704896540
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1704896540
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1704896540
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1704896540
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp 1704896540
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp 1704896540
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp 1704896540
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp 1704896540
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp 1704896540
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_63
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_66
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_68
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_69
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_72
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_89
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_92
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_93
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_95
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_96
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_98
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_99
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_101
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_102
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_104
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_105
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_107
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_108
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 1704896540
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_110
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_111
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 1704896540
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_113
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_114
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 1704896540
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_116
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_117
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 1704896540
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_119
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_120
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 1704896540
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_122
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_123
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 1704896540
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_125
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_126
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 1704896540
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_128
timestamp 1704896540
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_129
timestamp 1704896540
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 1704896540
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_131
timestamp 1704896540
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_132
timestamp 1704896540
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 1704896540
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_134
timestamp 1704896540
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_135
timestamp 1704896540
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 1704896540
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_137
timestamp 1704896540
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_138
timestamp 1704896540
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 1704896540
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_140
timestamp 1704896540
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_141
timestamp 1704896540
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 1704896540
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 1704896540
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 1704896540
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_145
timestamp 1704896540
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
<< labels >>
flabel metal4 s 2604 2128 2924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7604 2128 7924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12604 2128 12924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17604 2128 17924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3676 18908 3996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8676 18908 8996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 13676 18908 13996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6944 2128 7264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11944 2128 12264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 16944 2128 17264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3016 18908 3336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8016 18908 8336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 13016 18908 13336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 din1[0]
port 2 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 din1[1]
port 3 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 din1[2]
port 4 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 din1[3]
port 5 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 din1[4]
port 6 nsew signal input
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 din1[5]
port 7 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 din1[6]
port 8 nsew signal input
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 din1[7]
port 9 nsew signal input
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 din2[0]
port 10 nsew signal input
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 din2[1]
port 11 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 din2[2]
port 12 nsew signal input
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 din2[3]
port 13 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 din2[4]
port 14 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 din2[5]
port 15 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 din2[6]
port 16 nsew signal input
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 din2[7]
port 17 nsew signal input
flabel metal3 s 19200 18504 20000 18624 0 FreeSans 480 0 0 0 dout[0]
port 18 nsew signal output
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 dout[1]
port 19 nsew signal output
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 dout[2]
port 20 nsew signal output
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 dout[3]
port 21 nsew signal output
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 dout[4]
port 22 nsew signal output
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 dout[5]
port 23 nsew signal output
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 dout[6]
port 24 nsew signal output
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 480 0 0 0 dout[7]
port 25 nsew signal output
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 op[0]
port 26 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 op[1]
port 27 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 op[2]
port 28 nsew signal input
rlabel metal1 9982 17408 9982 17408 0 VGND
rlabel metal1 9982 16864 9982 16864 0 VPWR
rlabel metal1 2530 11084 2530 11084 0 _000_
rlabel metal1 9982 16728 9982 16728 0 _001_
rlabel metal2 15686 16898 15686 16898 0 _002_
rlabel metal1 2162 11220 2162 11220 0 _003_
rlabel metal1 8183 6426 8183 6426 0 _004_
rlabel metal1 14720 15470 14720 15470 0 _005_
rlabel metal2 4186 8840 4186 8840 0 _006_
rlabel via3 16859 12716 16859 12716 0 _007_
rlabel metal1 15962 13396 15962 13396 0 _008_
rlabel via3 6693 15300 6693 15300 0 _009_
rlabel metal2 17986 8993 17986 8993 0 _010_
rlabel metal2 7866 11713 7866 11713 0 _011_
rlabel metal1 15226 13362 15226 13362 0 _012_
rlabel via2 16146 2363 16146 2363 0 _013_
rlabel metal3 9223 2652 9223 2652 0 _014_
rlabel metal1 14812 13226 14812 13226 0 _015_
rlabel metal2 16146 6477 16146 6477 0 _016_
rlabel metal1 14582 14450 14582 14450 0 _017_
rlabel metal2 13202 16150 13202 16150 0 _018_
rlabel metal2 13018 13107 13018 13107 0 _019_
rlabel metal1 14076 15878 14076 15878 0 _020_
rlabel metal1 16330 8602 16330 8602 0 _021_
rlabel metal1 16744 2618 16744 2618 0 _022_
rlabel metal1 9016 14518 9016 14518 0 _023_
rlabel metal1 17572 2550 17572 2550 0 _024_
rlabel metal2 7590 14620 7590 14620 0 _025_
rlabel metal1 10534 11526 10534 11526 0 _026_
rlabel metal2 16514 8415 16514 8415 0 _027_
rlabel metal2 12558 6817 12558 6817 0 _028_
rlabel metal2 15410 4947 15410 4947 0 _029_
rlabel metal1 5382 13362 5382 13362 0 _030_
rlabel metal1 15272 5202 15272 5202 0 _031_
rlabel metal1 15824 5338 15824 5338 0 _032_
rlabel metal1 7544 14314 7544 14314 0 _033_
rlabel via3 15387 8228 15387 8228 0 _034_
rlabel via2 16882 15419 16882 15419 0 _035_
rlabel metal2 8326 14994 8326 14994 0 _036_
rlabel metal1 2484 8058 2484 8058 0 _037_
rlabel metal2 7636 8602 7636 8602 0 _038_
rlabel metal1 3956 7786 3956 7786 0 _039_
rlabel metal1 4600 8058 4600 8058 0 _040_
rlabel metal2 6026 10812 6026 10812 0 _041_
rlabel metal1 6072 15130 6072 15130 0 _042_
rlabel metal2 3634 5984 3634 5984 0 _043_
rlabel metal1 5842 3706 5842 3706 0 _044_
rlabel metal1 7222 8364 7222 8364 0 _045_
rlabel metal2 5750 9044 5750 9044 0 _046_
rlabel metal1 16422 5712 16422 5712 0 _047_
rlabel metal1 13202 12135 13202 12135 0 _048_
rlabel metal2 8418 15164 8418 15164 0 _049_
rlabel metal2 18262 6273 18262 6273 0 _050_
rlabel metal1 18216 6426 18216 6426 0 _051_
rlabel metal2 15410 11407 15410 11407 0 _052_
rlabel metal1 15134 3468 15134 3468 0 _053_
rlabel metal1 13110 5202 13110 5202 0 _054_
rlabel metal2 13018 11917 13018 11917 0 _055_
rlabel metal1 15088 3570 15088 3570 0 _056_
rlabel metal1 16330 3706 16330 3706 0 _057_
rlabel metal1 13754 15368 13754 15368 0 _058_
rlabel metal1 15364 12750 15364 12750 0 _059_
rlabel metal1 13018 12614 13018 12614 0 _060_
rlabel metal1 12604 10982 12604 10982 0 _061_
rlabel metal2 1518 10336 1518 10336 0 _062_
rlabel metal1 15640 7514 15640 7514 0 _063_
rlabel metal1 14168 4454 14168 4454 0 _064_
rlabel metal2 14122 5015 14122 5015 0 _065_
rlabel metal1 15916 10438 15916 10438 0 _066_
rlabel metal2 5566 9571 5566 9571 0 _067_
rlabel metal1 5658 4080 5658 4080 0 _068_
rlabel metal1 14168 15674 14168 15674 0 _069_
rlabel metal2 18124 15572 18124 15572 0 _070_
rlabel metal1 4922 10132 4922 10132 0 _071_
rlabel metal1 16008 16422 16008 16422 0 _072_
rlabel metal1 1518 2346 1518 2346 0 _073_
rlabel metal1 8280 7854 8280 7854 0 _074_
rlabel metal2 8326 7548 8326 7548 0 _075_
rlabel metal1 16836 4794 16836 4794 0 _076_
rlabel metal1 4922 2414 4922 2414 0 _077_
rlabel metal1 1610 2550 1610 2550 0 _078_
rlabel metal1 10534 6426 10534 6426 0 _079_
rlabel metal1 14306 16456 14306 16456 0 _080_
rlabel via1 12535 3026 12535 3026 0 _081_
rlabel via3 10971 15300 10971 15300 0 _082_
rlabel via2 1518 15963 1518 15963 0 _083_
rlabel metal1 16652 14790 16652 14790 0 _084_
rlabel metal2 7038 8636 7038 8636 0 _085_
rlabel metal1 12006 3060 12006 3060 0 _086_
rlabel metal2 8970 3434 8970 3434 0 _087_
rlabel metal1 10074 2618 10074 2618 0 _088_
rlabel metal2 14398 3689 14398 3689 0 _089_
rlabel metal2 13294 7055 13294 7055 0 _090_
rlabel metal1 6670 16524 6670 16524 0 _091_
rlabel metal1 7268 12682 7268 12682 0 _092_
rlabel metal1 14306 11220 14306 11220 0 _093_
rlabel via2 13202 5117 13202 5117 0 _094_
rlabel metal1 14582 11084 14582 11084 0 _095_
rlabel metal1 12466 11152 12466 11152 0 _096_
rlabel metal2 17710 7905 17710 7905 0 _097_
rlabel metal1 16698 5882 16698 5882 0 _098_
rlabel metal1 18032 4046 18032 4046 0 _099_
rlabel metal1 15364 15402 15364 15402 0 _100_
rlabel metal2 1426 6290 1426 6290 0 _101_
rlabel metal2 3082 16031 3082 16031 0 _102_
rlabel metal1 1840 10642 1840 10642 0 _103_
rlabel metal1 15962 4454 15962 4454 0 _104_
rlabel metal2 5382 10098 5382 10098 0 _105_
rlabel metal2 12466 7021 12466 7021 0 _106_
rlabel metal2 2530 16626 2530 16626 0 _107_
rlabel metal1 16698 15470 16698 15470 0 _108_
rlabel metal2 15226 10370 15226 10370 0 _109_
rlabel metal1 14674 5304 14674 5304 0 _110_
rlabel metal1 13478 12954 13478 12954 0 _111_
rlabel metal1 14398 12818 14398 12818 0 _112_
rlabel metal1 16008 17170 16008 17170 0 _113_
rlabel metal1 8234 12750 8234 12750 0 _114_
rlabel metal2 15226 16881 15226 16881 0 _115_
rlabel metal2 2346 6120 2346 6120 0 _116_
rlabel via2 13570 15555 13570 15555 0 _117_
rlabel metal1 18262 9418 18262 9418 0 _118_
rlabel metal1 13570 13294 13570 13294 0 _119_
rlabel metal2 17066 14093 17066 14093 0 _120_
rlabel metal1 17158 14348 17158 14348 0 _121_
rlabel metal2 4002 14127 4002 14127 0 _122_
rlabel via2 14398 14909 14398 14909 0 _123_
rlabel metal1 16054 14382 16054 14382 0 _124_
rlabel metal1 13570 13362 13570 13362 0 _125_
rlabel metal2 13754 6409 13754 6409 0 _126_
rlabel metal1 13938 5882 13938 5882 0 _127_
rlabel metal1 18400 15402 18400 15402 0 _128_
rlabel metal1 15916 8466 15916 8466 0 _129_
rlabel metal1 15042 8908 15042 8908 0 _130_
rlabel metal2 14766 11866 14766 11866 0 _131_
rlabel metal1 14536 8806 14536 8806 0 _132_
rlabel metal1 14582 4590 14582 4590 0 _133_
rlabel metal1 1702 2448 1702 2448 0 _134_
rlabel metal1 12650 16490 12650 16490 0 _135_
rlabel metal1 13570 6222 13570 6222 0 _136_
rlabel metal1 9522 15538 9522 15538 0 _137_
rlabel metal1 13938 7174 13938 7174 0 _138_
rlabel metal3 13593 13804 13593 13804 0 _139_
rlabel via2 1794 6171 1794 6171 0 _140_
rlabel metal1 5566 12818 5566 12818 0 _141_
rlabel metal1 17342 15572 17342 15572 0 _142_
rlabel metal1 14168 13906 14168 13906 0 _143_
rlabel metal1 16054 13702 16054 13702 0 _144_
rlabel metal1 18032 15470 18032 15470 0 _145_
rlabel metal1 13654 7514 13654 7514 0 _146_
rlabel metal1 2162 2992 2162 2992 0 _147_
rlabel metal1 2553 3026 2553 3026 0 _148_
rlabel metal3 16767 15572 16767 15572 0 _149_
rlabel metal1 18216 16082 18216 16082 0 _150_
rlabel metal2 15502 15844 15502 15844 0 _151_
rlabel metal2 3174 4709 3174 4709 0 _152_
rlabel metal1 15226 4998 15226 4998 0 _153_
rlabel metal1 18308 16694 18308 16694 0 _154_
rlabel metal1 10442 12784 10442 12784 0 _155_
rlabel metal2 14214 7650 14214 7650 0 _156_
rlabel metal1 8372 13974 8372 13974 0 _157_
rlabel metal2 13478 4420 13478 4420 0 _158_
rlabel metal1 2346 9486 2346 9486 0 _159_
rlabel metal4 2484 6732 2484 6732 0 _160_
rlabel metal1 16652 16558 16652 16558 0 _161_
rlabel metal2 14674 16796 14674 16796 0 _162_
rlabel metal1 9384 6970 9384 6970 0 _163_
rlabel metal1 8510 13498 8510 13498 0 _164_
rlabel metal2 15778 2465 15778 2465 0 _165_
rlabel metal1 14306 8602 14306 8602 0 _166_
rlabel via2 14214 16507 14214 16507 0 _167_
rlabel metal1 7222 6630 7222 6630 0 _168_
rlabel metal2 15594 13532 15594 13532 0 _169_
rlabel metal3 751 9316 751 9316 0 din1[0]
rlabel metal3 1050 8228 1050 8228 0 din1[1]
rlabel metal3 751 7140 751 7140 0 din1[2]
rlabel metal3 820 6052 820 6052 0 din1[3]
rlabel metal3 751 4964 751 4964 0 din1[4]
rlabel metal3 751 3876 751 3876 0 din1[5]
rlabel metal3 751 2788 751 2788 0 din1[6]
rlabel metal3 1280 1700 1280 1700 0 din1[7]
rlabel metal3 1280 18020 1280 18020 0 din2[0]
rlabel metal3 751 16932 751 16932 0 din2[1]
rlabel metal3 866 15844 866 15844 0 din2[2]
rlabel metal3 751 14756 751 14756 0 din2[3]
rlabel metal3 1050 13668 1050 13668 0 din2[4]
rlabel metal3 751 12580 751 12580 0 din2[5]
rlabel metal3 751 11492 751 11492 0 din2[6]
rlabel metal3 751 10404 751 10404 0 din2[7]
rlabel metal1 18216 17306 18216 17306 0 dout[0]
rlabel metal1 17664 16422 17664 16422 0 dout[1]
rlabel metal2 18446 13855 18446 13855 0 dout[2]
rlabel metal2 18446 11373 18446 11373 0 dout[3]
rlabel via2 18446 8789 18446 8789 0 dout[4]
rlabel metal2 18446 6477 18446 6477 0 dout[5]
rlabel via2 18446 3893 18446 3893 0 dout[6]
rlabel metal2 18446 1853 18446 1853 0 dout[7]
rlabel metal1 1610 9656 1610 9656 0 net1
rlabel metal1 10028 12138 10028 12138 0 net10
rlabel metal1 9292 6698 9292 6698 0 net11
rlabel metal2 15134 10404 15134 10404 0 net12
rlabel metal1 1702 13702 1702 13702 0 net13
rlabel metal1 1748 12954 1748 12954 0 net14
rlabel metal1 2898 7854 2898 7854 0 net15
rlabel metal1 8004 5134 8004 5134 0 net16
rlabel metal2 9430 14994 9430 14994 0 net17
rlabel metal1 12880 2550 12880 2550 0 net18
rlabel metal1 4416 2618 4416 2618 0 net19
rlabel metal1 12834 5236 12834 5236 0 net2
rlabel metal2 18262 17340 18262 17340 0 net20
rlabel via2 5106 10149 5106 10149 0 net21
rlabel metal1 16790 13906 16790 13906 0 net22
rlabel metal1 15686 2822 15686 2822 0 net23
rlabel metal1 17710 8058 17710 8058 0 net24
rlabel metal1 17940 16626 17940 16626 0 net25
rlabel metal2 18262 4862 18262 4862 0 net26
rlabel metal1 18446 2414 18446 2414 0 net27
rlabel metal1 11960 4590 11960 4590 0 net28
rlabel metal1 1748 7446 1748 7446 0 net3
rlabel metal2 13018 14875 13018 14875 0 net4
rlabel metal1 2070 9996 2070 9996 0 net5
rlabel metal1 12512 13974 12512 13974 0 net6
rlabel metal2 1702 5134 1702 5134 0 net7
rlabel metal1 13892 5678 13892 5678 0 net8
rlabel metal1 1702 16966 1702 16966 0 net9
rlabel metal2 16606 1588 16606 1588 0 op[0]
rlabel metal2 9982 1554 9982 1554 0 op[1]
rlabel metal2 3358 1554 3358 1554 0 op[2]
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
